--------------------------------------------------------------------------------
--
-- File Type:    VHDL 
-- Tool Version: verilog2vhdl 19.00c
-- Input file was: ./netlists/module_fnChkNodeCore.vg.vpp
-- Command line was: /home/sandeep/Desktop/ActualCoursework/SemII/EE705/synapticad-19.00c-x64/bin/x86_64/verilog2vhdl.bin ./netlists/module_fnChkNodeCore.vg -No_Component_Check
-- Date Created: Sat Apr 27 19:23:32 2019
--
--------------------------------------------------------------------------------



LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY ASC;
USE ASC.numeric_std.all;
ENTITY module_fnChkNodeCore IS	-- 
    PORT (
        SIGNAL fnChkNodeCore_i_0 : IN std_logic;	
        SIGNAL fnChkNodeCore_i_1 : IN std_logic;	
        SIGNAL fnChkNodeCore_i_2 : IN std_logic;	
        SIGNAL fnChkNodeCore_0 : OUT std_logic;	
        SIGNAL fnChkNodeCore_1 : OUT std_logic;	
        SIGNAL fnChkNodeCore_2 : OUT std_logic);	
END module_fnChkNodeCore;

-- /* Generated by Yosys 0.7 (git sha1 61f6811, gcc 5.4.0-6ubuntu1~16.04.4 -O2 -fstack-protector-strong -fPIC -Os) */

LIBRARY ASC;

LIBRARY user_defined;
ARCHITECTURE VeriArch OF module_fnChkNodeCore IS
    USE ASC.FUNCTIONS.ALL;
    USE user_defined.user_package.ALL;

    SIGNAL ag_00 : std_logic;	

    SIGNAL ag_01 : std_logic;	

    SIGNAL ag_02 : std_logic;	

    SIGNAL ag_03 : std_logic;	

    SIGNAL ag_04 : std_logic;	

    SIGNAL ag_05 : std_logic;	

    SIGNAL ag_06 : std_logic;	

    SIGNAL ag_07 : std_logic;	

    SIGNAL ag_08 : std_logic;	
-- Intermediate signal for fnChkNodeCore_0
    SIGNAL V2V_fnChkNodeCore_0 : std_logic;	
-- Intermediate signal for fnChkNodeCore_1
    SIGNAL V2V_fnChkNodeCore_1 : std_logic;	
-- Intermediate signal for fnChkNodeCore_2
    SIGNAL V2V_fnChkNodeCore_2 : std_logic;	

    SIGNAL GUARD : boolean:= TRUE;	
BEGIN
    fnChkNodeCore_0 <= V2V_fnChkNodeCore_0;	
    fnChkNodeCore_1 <= V2V_fnChkNodeCore_1;	
    fnChkNodeCore_2 <= V2V_fnChkNodeCore_2;	

    ag_09 : user_defined.user_package.std_inv
    PORT MAP (
        a => fnChkNodeCore_i_2,
        y => ag_06);	


    ag_10 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_06,
        b => fnChkNodeCore_i_1,
        y => ag_07);	


    ag_11 : user_defined.user_package.std_inv
    PORT MAP (
        a => fnChkNodeCore_i_1,
        y => ag_08);	


    ag_12 : user_defined.user_package.std_nand2
    PORT MAP (
        a => fnChkNodeCore_i_2,
        b => ag_08,
        y => ag_00);	


    ag_13 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_00,
        b => ag_07,
        y => V2V_fnChkNodeCore_0);	


    ag_14 : user_defined.user_package.std_inv
    PORT MAP (
        a => fnChkNodeCore_i_0,
        y => ag_01);	


    ag_15 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_01,
        b => fnChkNodeCore_i_2,
        y => ag_02);	


    ag_16 : user_defined.user_package.std_nand2
    PORT MAP (
        a => fnChkNodeCore_i_0,
        b => ag_06,
        y => ag_03);	


    ag_17 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_03,
        b => ag_02,
        y => V2V_fnChkNodeCore_1);	


    ag_18 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_01,
        b => fnChkNodeCore_i_1,
        y => ag_04);	


    ag_19 : user_defined.user_package.std_nand2
    PORT MAP (
        a => fnChkNodeCore_i_0,
        b => ag_08,
        y => ag_05);	


    ag_20 : user_defined.user_package.std_nand2
    PORT MAP (
        a => ag_05,
        b => ag_04,
        y => V2V_fnChkNodeCore_2);	

END VeriArch;

