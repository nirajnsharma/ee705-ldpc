module std_inv(a,y);
input a;
output y;
assign y=~a;
endmodule