--------------------------------------------------------------------------------
--
-- File Type:    VHDL 
-- Tool Version: verilog2vhdl 19.00c
-- Input file was: ./module_fnBitNodeCore.vg.vpp
-- Command line was: /home/sandeep/Desktop/ActualCoursework/SemII/EE705/synapticad-19.00c-x64/bin/x86_64/verilog2vhdl.bin ./module_fnBitNodeCore.vg -No_Component_Check
-- Date Created: Sat Apr 27 18:28:47 2019
--
--------------------------------------------------------------------------------



LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY ASC;
USE ASC.numeric_std.all;
ENTITY module_fnBitNodeCore IS	-- 
    PORT (
        SIGNAL \fnBitNodeCore_i[0]\ : IN std_logic;	
        SIGNAL \fnBitNodeCore_i[1]\ : IN std_logic;	
        SIGNAL \fnBitNodeCore_i[2]\ : IN std_logic;	
        SIGNAL fnBitNodeCore : OUT std_logic);	
END module_fnBitNodeCore;

-- /* Generated by Yosys 0.7 (git sha1 61f6811, gcc 5.4.0-6ubuntu1~16.04.4 -O2 -fstack-protector-strong -fPIC -Os) */

LIBRARY ASC;

LIBRARY user_defined;
ARCHITECTURE VeriArch OF module_fnBitNodeCore IS
    USE ASC.FUNCTIONS.ALL;
    USE user_defined.user_package.ALL;

    SIGNAL \ag_00_\ : std_logic;	

    SIGNAL \ag_01_\ : std_logic;	

    SIGNAL \ag_02_\ : std_logic;	

    SIGNAL \ag_03_\ : std_logic;	

    SIGNAL \ag_04_\ : std_logic;	
-- Intermediate signal for fnBitNodeCore
    SIGNAL V2V_fnBitNodeCore : std_logic;	

    SIGNAL GUARD : boolean:= TRUE;	
BEGIN
    fnBitNodeCore <= V2V_fnBitNodeCore;	

    \ag_05_\ : user_defined.user_package.std_nand2
    PORT MAP (
        a => \fnBitNodeCore_i[0]\,
        b => \fnBitNodeCore_i[1]\,
        y => \ag_00_\);	


    \ag_06_\ : user_defined.user_package.std_inv
    PORT MAP (
        a => \fnBitNodeCore_i[1]\,
        y => \ag_01_\);	


    \ag_07_\ : user_defined.user_package.std_inv
    PORT MAP (
        a => \fnBitNodeCore_i[0]\,
        y => \ag_02_\);	


    \ag_08_\ : user_defined.user_package.std_nand2
    PORT MAP (
        a => \ag_02_\,
        b => \ag_01_\,
        y => \ag_03_\);	


    \ag_09_\ : user_defined.user_package.std_nand2
    PORT MAP (
        a => \ag_03_\,
        b => \fnBitNodeCore_i[2]\,
        y => \ag_04_\);	


    \ag_10_\ : user_defined.user_package.std_nand2
    PORT MAP (
        a => \ag_04_\,
        b => \ag_00_\,
        y => V2V_fnBitNodeCore);	

END VeriArch;

