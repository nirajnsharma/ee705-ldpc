magic
tech scmos
magscale 1 2
timestamp 1556798218
<< metal1 >>
rect 3272 5806 3278 5814
rect 3286 5806 3292 5814
rect 3300 5806 3306 5814
rect 3314 5806 3320 5814
rect 6344 5806 6350 5814
rect 6358 5806 6364 5814
rect 6372 5806 6378 5814
rect 6386 5806 6392 5814
rect 948 5756 956 5764
rect 1492 5757 1524 5763
rect 1516 5748 1524 5757
rect 1868 5752 1876 5756
rect 253 5737 275 5743
rect 349 5737 364 5743
rect 653 5737 675 5743
rect 893 5737 947 5743
rect 1320 5736 1324 5744
rect 1677 5737 1692 5743
rect 2429 5737 2451 5743
rect 2749 5737 2771 5743
rect 3165 5737 3187 5743
rect 3693 5737 3715 5743
rect 4125 5737 4147 5743
rect 5508 5737 5523 5743
rect 5620 5737 5635 5743
rect 6109 5737 6131 5743
rect 7037 5737 7052 5743
rect 77 5717 92 5723
rect 212 5717 227 5723
rect 1044 5717 1059 5723
rect 1181 5717 1219 5723
rect 1213 5697 1219 5717
rect 1661 5717 1676 5723
rect 1709 5717 1788 5723
rect 2253 5717 2268 5723
rect 2292 5717 2307 5723
rect 2388 5717 2403 5723
rect 2509 5723 2515 5736
rect 2509 5717 2531 5723
rect 2717 5717 2732 5723
rect 2797 5717 2812 5723
rect 2932 5717 2947 5723
rect 3133 5717 3148 5723
rect 3213 5717 3276 5723
rect 3805 5723 3811 5736
rect 3757 5717 3795 5723
rect 3805 5717 3827 5723
rect 1284 5697 1299 5703
rect 3757 5697 3763 5717
rect 4029 5723 4035 5736
rect 4013 5717 4035 5723
rect 4045 5717 4083 5723
rect 4077 5697 4083 5717
rect 5101 5717 5155 5723
rect 5405 5717 5443 5723
rect 5501 5717 5523 5723
rect 5549 5717 5612 5723
rect 5517 5704 5523 5717
rect 5645 5717 5667 5723
rect 5988 5716 5992 5724
rect 7069 5717 7100 5723
rect 7268 5696 7272 5704
rect 621 5677 636 5683
rect 1242 5676 1244 5684
rect 1510 5676 1516 5684
rect 4212 5676 4218 5684
rect 5334 5676 5340 5684
rect 1818 5636 1820 5644
rect 7400 5636 7404 5644
rect 1736 5606 1742 5614
rect 1750 5606 1756 5614
rect 1764 5606 1770 5614
rect 1778 5606 1784 5614
rect 4808 5606 4814 5614
rect 4822 5606 4828 5614
rect 4836 5606 4842 5614
rect 4850 5606 4856 5614
rect 362 5576 364 5584
rect 2250 5576 2252 5584
rect 2340 5576 2342 5584
rect 4116 5576 4118 5584
rect 4500 5576 4502 5584
rect 6004 5576 6006 5584
rect 6756 5576 6758 5584
rect 7284 5576 7286 5584
rect 1930 5556 1932 5564
rect 4378 5556 4380 5564
rect 4810 5556 4812 5564
rect 5908 5556 5910 5564
rect 7946 5556 7948 5564
rect 500 5537 515 5543
rect 2036 5537 2051 5543
rect 2156 5537 2172 5543
rect 5028 5537 5043 5543
rect 5098 5536 5100 5544
rect 5780 5536 5782 5544
rect 7092 5537 7107 5543
rect 7348 5537 7363 5543
rect 8004 5536 8006 5544
rect 436 5497 467 5503
rect 637 5497 659 5503
rect 1085 5503 1091 5523
rect 1060 5497 1075 5503
rect 1085 5497 1123 5503
rect 1325 5497 1356 5503
rect 1469 5503 1475 5523
rect 1885 5517 1907 5523
rect 2045 5517 2067 5523
rect 2653 5517 2691 5523
rect 4301 5517 4332 5523
rect 4964 5516 4972 5524
rect 5933 5517 5971 5523
rect 6077 5517 6099 5523
rect 7309 5517 7331 5523
rect 8029 5517 8067 5523
rect 1469 5497 1507 5503
rect 1517 5497 1539 5503
rect 1668 5497 1683 5503
rect 2100 5497 2131 5503
rect 2141 5497 2156 5503
rect 2189 5497 2220 5503
rect 2349 5497 2371 5503
rect 2772 5497 2787 5503
rect 2925 5497 2940 5503
rect 3309 5497 3324 5503
rect 3444 5497 3459 5503
rect 4052 5497 4067 5503
rect 4141 5497 4179 5503
rect 4452 5497 4483 5503
rect 429 5477 451 5483
rect 445 5464 451 5477
rect 612 5477 627 5483
rect 1348 5477 1363 5483
rect 2269 5477 2291 5483
rect 2733 5477 2755 5483
rect 3181 5477 3212 5483
rect 3485 5477 3507 5483
rect 4477 5477 4483 5497
rect 4765 5497 4780 5503
rect 4813 5497 4915 5503
rect 5053 5497 5068 5503
rect 5764 5497 5779 5503
rect 6036 5497 6067 5503
rect 6157 5497 6179 5503
rect 6196 5497 6212 5503
rect 6204 5492 6212 5497
rect 6333 5497 6419 5503
rect 5965 5477 5987 5483
rect 6333 5483 6339 5497
rect 6644 5497 6659 5503
rect 6669 5497 6684 5503
rect 6836 5497 6851 5503
rect 7197 5497 7219 5503
rect 7565 5497 7587 5503
rect 8061 5497 8076 5503
rect 6301 5477 6339 5483
rect 6605 5477 6620 5483
rect 6717 5477 6739 5483
rect 2388 5457 2403 5463
rect 4132 5457 4147 5463
rect 4157 5457 4172 5463
rect 5220 5457 5235 5463
rect 1741 5437 1756 5443
rect 2826 5436 2828 5444
rect 3162 5436 3164 5444
rect 4234 5436 4236 5444
rect 3272 5406 3278 5414
rect 3286 5406 3292 5414
rect 3300 5406 3306 5414
rect 3314 5406 3320 5414
rect 6344 5406 6350 5414
rect 6358 5406 6364 5414
rect 6372 5406 6378 5414
rect 6386 5406 6392 5414
rect 1844 5376 1848 5384
rect 3626 5376 3628 5384
rect 6554 5376 6556 5384
rect 7908 5377 7923 5383
rect 765 5357 787 5363
rect 2013 5357 2028 5363
rect 4973 5357 4988 5363
rect 5204 5356 5212 5364
rect 5309 5357 5347 5363
rect 5357 5357 5372 5363
rect 5524 5357 5539 5363
rect 6605 5357 6620 5363
rect 605 5337 620 5343
rect 1325 5337 1347 5343
rect 1741 5337 1811 5343
rect 3149 5337 3164 5343
rect 3965 5337 4003 5343
rect 4077 5337 4108 5343
rect 468 5317 499 5323
rect 685 5317 739 5323
rect 852 5317 883 5323
rect 1508 5317 1523 5323
rect 1629 5317 1667 5323
rect 2036 5317 2051 5323
rect 2285 5317 2323 5323
rect 500 5296 508 5304
rect 589 5297 611 5303
rect 1277 5297 1292 5303
rect 2317 5297 2323 5317
rect 3133 5317 3180 5323
rect 3828 5317 3843 5323
rect 4020 5317 4035 5323
rect 4077 5317 4083 5337
rect 4292 5337 4307 5343
rect 5037 5337 5091 5343
rect 6285 5337 6307 5343
rect 6365 5337 6380 5343
rect 6653 5343 6659 5356
rect 6653 5337 6675 5343
rect 8036 5337 8051 5343
rect 5325 5317 5340 5323
rect 5373 5317 5395 5323
rect 5917 5317 5939 5323
rect 6084 5317 6099 5323
rect 6324 5317 6355 5323
rect 7188 5317 7203 5323
rect 3020 5303 3028 5308
rect 3020 5297 3043 5303
rect 6228 5297 6243 5303
rect 6509 5297 6547 5303
rect 7028 5296 7036 5304
rect 7053 5297 7068 5303
rect 7197 5297 7203 5317
rect 7277 5317 7292 5323
rect 7460 5317 7475 5323
rect 8052 5317 8083 5323
rect 7293 5297 7315 5303
rect 7780 5297 7795 5303
rect 7292 5284 7300 5288
rect 564 5276 566 5284
rect 2790 5276 2796 5284
rect 4365 5277 4419 5283
rect 7444 5256 7446 5264
rect 1620 5236 1622 5244
rect 7850 5236 7852 5244
rect 1736 5206 1742 5214
rect 1750 5206 1756 5214
rect 1764 5206 1770 5214
rect 1778 5206 1784 5214
rect 4808 5206 4814 5214
rect 4822 5206 4828 5214
rect 4836 5206 4842 5214
rect 4850 5206 4856 5214
rect 1789 5177 1804 5183
rect 6180 5176 6182 5184
rect 7780 5176 7782 5184
rect 6244 5156 6246 5164
rect 540 5132 548 5136
rect 2340 5136 2344 5144
rect 2524 5137 2540 5143
rect 3786 5136 3788 5144
rect 7101 5137 7116 5143
rect 7613 5137 7628 5143
rect 668 5132 676 5136
rect 4828 5132 4836 5136
rect 276 5097 307 5103
rect 413 5097 435 5103
rect 621 5097 659 5103
rect 861 5097 876 5103
rect 1524 5097 1539 5103
rect 2125 5103 2131 5123
rect 2413 5117 2444 5123
rect 2061 5097 2083 5103
rect 2093 5097 2131 5103
rect 2909 5103 2915 5123
rect 2964 5117 2979 5123
rect 2909 5097 2947 5103
rect 3268 5097 3331 5103
rect 3517 5103 3523 5123
rect 3501 5097 3523 5103
rect 3668 5097 3683 5103
rect 3892 5097 3923 5103
rect 4381 5097 4403 5103
rect 4564 5097 4579 5103
rect 4884 5097 4899 5103
rect 4957 5097 4995 5103
rect 5053 5097 5068 5103
rect 5220 5097 5235 5103
rect 5325 5097 5347 5103
rect 5485 5097 5507 5103
rect 7085 5103 7091 5123
rect 7684 5116 7692 5124
rect 7981 5117 7996 5123
rect 6973 5097 6995 5103
rect 7053 5097 7091 5103
rect 7373 5097 7395 5103
rect 7956 5097 7971 5103
rect 7340 5092 7348 5096
rect 1400 5076 1404 5084
rect 2244 5077 2275 5083
rect 2285 5077 2300 5083
rect 2461 5077 2476 5083
rect 2637 5077 2659 5083
rect 3245 5077 3315 5083
rect 3485 5077 3500 5083
rect 3661 5077 3676 5083
rect 3805 5077 3827 5083
rect 4669 5077 4691 5083
rect 4756 5077 4771 5083
rect 5069 5077 5091 5083
rect 5260 5066 5268 5076
rect 5421 5077 5436 5083
rect 1165 5057 1187 5063
rect 3588 5057 3603 5063
rect 1268 5036 1270 5044
rect 2900 5036 2902 5044
rect 3866 5036 3868 5044
rect 4349 5037 4355 5063
rect 4420 5057 4435 5063
rect 5373 5057 5395 5063
rect 5421 5057 5427 5077
rect 5885 5077 5907 5083
rect 6068 5076 6070 5084
rect 6445 5077 6460 5083
rect 7181 5077 7203 5083
rect 7645 5077 7667 5083
rect 7741 5077 7763 5083
rect 7837 5077 7891 5083
rect 7940 5077 7955 5083
rect 4829 5037 4876 5043
rect 5389 5037 5395 5057
rect 7396 5057 7411 5063
rect 5725 5037 5740 5043
rect 5810 5037 5836 5043
rect 3272 5006 3278 5014
rect 3286 5006 3292 5014
rect 3300 5006 3306 5014
rect 3314 5006 3320 5014
rect 6344 5006 6350 5014
rect 6358 5006 6364 5014
rect 6372 5006 6378 5014
rect 6386 5006 6392 5014
rect 1064 4976 1068 4984
rect 1220 4976 1222 4984
rect 3268 4976 3270 4984
rect 3444 4976 3446 4984
rect 5514 4976 5516 4984
rect 8074 4976 8076 4984
rect 4724 4956 4732 4964
rect 420 4937 440 4943
rect 477 4937 499 4943
rect 1101 4937 1123 4943
rect 1236 4937 1251 4943
rect 2484 4937 2499 4943
rect 2621 4937 2636 4943
rect 2877 4937 2899 4943
rect 3197 4937 3219 4943
rect 3236 4937 3251 4943
rect 3284 4937 3347 4943
rect 3853 4937 3875 4943
rect 4413 4937 4435 4943
rect 4637 4937 4659 4943
rect 5629 4943 5635 4963
rect 5836 4957 5868 4963
rect 5836 4948 5844 4957
rect 6220 4957 6243 4963
rect 6220 4954 6228 4957
rect 5597 4937 5619 4943
rect 5629 4937 5644 4943
rect 5661 4937 5699 4943
rect 6253 4937 6275 4943
rect 6340 4937 6387 4943
rect 6717 4937 6748 4943
rect 6904 4937 6924 4943
rect 61 4917 115 4923
rect 253 4917 268 4923
rect 525 4917 556 4923
rect 573 4917 604 4923
rect 1165 4917 1196 4923
rect 1341 4917 1379 4923
rect 1405 4917 1443 4923
rect 244 4896 252 4904
rect 628 4896 636 4904
rect 1373 4897 1379 4917
rect 1565 4917 1603 4923
rect 2541 4917 2572 4923
rect 2861 4917 2876 4923
rect 3156 4917 3171 4923
rect 3453 4917 3491 4923
rect 2205 4897 2220 4903
rect 2852 4896 2860 4904
rect 3277 4897 3292 4903
rect 3300 4897 3340 4903
rect 3373 4897 3388 4903
rect 3453 4897 3459 4917
rect 3837 4917 3852 4923
rect 4237 4917 4252 4923
rect 4372 4917 4387 4923
rect 4397 4917 4412 4923
rect 6548 4917 6563 4923
rect 6653 4917 6668 4923
rect 6804 4917 6835 4923
rect 7684 4917 7699 4923
rect 7780 4917 7795 4923
rect 7869 4917 7923 4923
rect 8029 4917 8067 4923
rect 6588 4904 6596 4914
rect 5677 4897 5692 4903
rect 5764 4896 5772 4904
rect 6932 4897 6947 4903
rect 7700 4896 7708 4904
rect 7757 4897 7772 4903
rect 8061 4897 8067 4917
rect 4716 4884 4724 4888
rect 5500 4884 5508 4888
rect 540 4877 556 4883
rect 2086 4876 2092 4884
rect 2148 4877 2163 4883
rect 2157 4857 2163 4877
rect 3405 4877 3420 4883
rect 4804 4877 4819 4883
rect 5996 4884 6004 4888
rect 5788 4877 5811 4883
rect 8100 4877 8131 4883
rect 1268 4836 1270 4844
rect 7866 4836 7868 4844
rect 1736 4806 1742 4814
rect 1750 4806 1756 4814
rect 1764 4806 1770 4814
rect 1778 4806 1784 4814
rect 4808 4806 4814 4814
rect 4822 4806 4828 4814
rect 4836 4806 4842 4814
rect 4850 4806 4856 4814
rect 5556 4776 5558 4784
rect 6996 4776 6998 4784
rect 5114 4756 5116 4764
rect 1828 4737 1843 4743
rect 2132 4736 2134 4744
rect 2596 4737 2611 4743
rect 2826 4736 2828 4744
rect 3780 4736 3782 4744
rect 5272 4736 5276 4744
rect 5972 4737 5987 4743
rect 7892 4737 7907 4743
rect 621 4717 652 4723
rect 1133 4697 1155 4703
rect 1533 4703 1539 4723
rect 2477 4717 2499 4723
rect 1421 4697 1475 4703
rect 1533 4697 1571 4703
rect 1757 4697 1779 4703
rect 221 4677 243 4683
rect 717 4677 771 4683
rect 797 4677 812 4683
rect 1757 4683 1763 4697
rect 2116 4697 2131 4703
rect 2189 4697 2227 4703
rect 2333 4697 2364 4703
rect 2532 4697 2563 4703
rect 2573 4697 2588 4703
rect 3613 4697 3667 4703
rect 3805 4703 3811 4723
rect 3805 4697 3843 4703
rect 3853 4697 3891 4703
rect 4020 4697 4051 4703
rect 4637 4703 4643 4723
rect 4868 4717 4883 4723
rect 4621 4697 4643 4703
rect 4692 4697 4723 4703
rect 4813 4697 4828 4703
rect 5004 4703 5012 4708
rect 5004 4697 5027 4703
rect 1613 4677 1667 4683
rect 1693 4677 1763 4683
rect 1860 4677 1875 4683
rect 2205 4677 2220 4683
rect 2269 4677 2323 4683
rect 4541 4677 4556 4683
rect 4628 4677 4643 4683
rect 4797 4677 4899 4683
rect 4972 4677 4988 4683
rect 4972 4676 4980 4677
rect 5021 4677 5027 4697
rect 5085 4703 5091 4723
rect 5053 4697 5091 4703
rect 5421 4697 5475 4703
rect 5581 4703 5587 4723
rect 5581 4697 5619 4703
rect 5837 4697 5852 4703
rect 5940 4697 5955 4703
rect 6637 4703 6643 4723
rect 6637 4697 6675 4703
rect 6941 4697 6956 4703
rect 7101 4703 7107 4723
rect 7444 4716 7452 4724
rect 7076 4697 7107 4703
rect 7165 4697 7187 4703
rect 7469 4703 7475 4723
rect 7677 4717 7692 4723
rect 8068 4716 8072 4724
rect 7469 4697 7507 4703
rect 7613 4697 7628 4703
rect 7812 4697 7827 4703
rect 7933 4697 7948 4703
rect 6028 4692 6036 4696
rect 5309 4677 5324 4683
rect 5885 4677 5907 4683
rect 6125 4677 6140 4683
rect 5885 4664 5891 4677
rect 7620 4677 7651 4683
rect 324 4656 332 4664
rect 1524 4656 1532 4664
rect 2500 4656 2508 4664
rect 5373 4657 5395 4663
rect 5965 4657 5987 4663
rect 6349 4657 6396 4663
rect 6804 4657 6819 4663
rect 6836 4657 6851 4663
rect 7108 4656 7116 4664
rect 7860 4656 7868 4664
rect 5924 4636 5926 4644
rect 6106 4636 6108 4644
rect 6372 4637 6419 4643
rect 6628 4636 6630 4644
rect 7572 4636 7574 4644
rect 3272 4606 3278 4614
rect 3286 4606 3292 4614
rect 3300 4606 3306 4614
rect 3314 4606 3320 4614
rect 6344 4606 6350 4614
rect 6358 4606 6364 4614
rect 6372 4606 6378 4614
rect 6386 4606 6392 4614
rect 3496 4576 3500 4584
rect 4660 4576 4662 4584
rect 7572 4576 7574 4584
rect 285 4557 300 4563
rect 541 4557 563 4563
rect 877 4557 899 4563
rect 1748 4557 1780 4563
rect 349 4543 355 4556
rect 1772 4548 1780 4557
rect 3332 4557 3363 4563
rect 349 4537 371 4543
rect 504 4536 508 4544
rect 941 4537 979 4543
rect 1620 4537 1636 4543
rect 2605 4537 2627 4543
rect 3428 4537 3443 4543
rect 3805 4537 3820 4543
rect 4100 4537 4147 4543
rect 4285 4537 4307 4543
rect 5677 4537 5715 4543
rect 5741 4537 5756 4543
rect 6548 4537 6563 4543
rect 6717 4537 6739 4543
rect 6772 4537 6812 4543
rect 6845 4537 6899 4543
rect 7588 4537 7603 4543
rect 7613 4537 7644 4543
rect 204 4524 212 4528
rect 100 4517 131 4523
rect 333 4517 364 4523
rect 564 4517 579 4523
rect 589 4517 611 4523
rect 925 4517 940 4523
rect 1276 4524 1284 4528
rect 2676 4517 2707 4523
rect 3373 4517 3395 4523
rect 3549 4517 3580 4523
rect 3885 4517 3916 4523
rect 4036 4517 4051 4523
rect 4196 4517 4211 4523
rect 4669 4517 4707 4523
rect 2573 4497 2611 4503
rect 2724 4497 2739 4503
rect 3293 4497 3308 4503
rect 3684 4497 3699 4503
rect 4228 4497 4243 4503
rect 4564 4496 4568 4504
rect 4669 4497 4675 4517
rect 5149 4517 5203 4523
rect 5229 4517 5267 4523
rect 5277 4517 5299 4523
rect 5229 4497 5235 4517
rect 5428 4517 5443 4523
rect 5572 4517 5603 4523
rect 5620 4517 5651 4523
rect 5661 4517 5676 4523
rect 5892 4517 5907 4523
rect 6141 4517 6195 4523
rect 6541 4517 6563 4523
rect 6589 4517 6604 4523
rect 6557 4504 6563 4517
rect 7405 4517 7459 4523
rect 7629 4517 7667 4523
rect 7629 4497 7635 4517
rect 7860 4517 7875 4523
rect 285 4477 300 4483
rect 452 4476 454 4484
rect 1380 4476 1386 4484
rect 2420 4476 2422 4484
rect 2548 4476 2550 4484
rect 2916 4476 2920 4484
rect 3126 4476 3132 4484
rect 3956 4477 3987 4483
rect 3981 4457 3987 4477
rect 4884 4476 4890 4484
rect 7796 4476 7802 4484
rect 1844 4437 1875 4443
rect 4052 4436 4054 4444
rect 1736 4406 1742 4414
rect 1750 4406 1756 4414
rect 1764 4406 1770 4414
rect 1778 4406 1784 4414
rect 4808 4406 4814 4414
rect 4822 4406 4828 4414
rect 4836 4406 4842 4414
rect 4850 4406 4856 4414
rect 868 4376 872 4384
rect 1082 4376 1084 4384
rect 1476 4376 1478 4384
rect 2804 4376 2806 4384
rect 3316 4377 3363 4383
rect 7626 4356 7628 4364
rect 948 4337 963 4343
rect 1901 4337 1924 4343
rect 2061 4337 2076 4343
rect 2212 4336 2214 4344
rect 2276 4336 2278 4344
rect 2698 4336 2700 4344
rect 3373 4337 3452 4343
rect 4468 4337 4483 4343
rect 4925 4337 4940 4343
rect 5716 4336 5718 4344
rect 6074 4336 6076 4344
rect 6756 4336 6760 4344
rect 7780 4337 7796 4343
rect 8092 4332 8100 4336
rect 4396 4324 4404 4328
rect 93 4303 99 4323
rect 740 4317 755 4323
rect 1012 4316 1020 4324
rect 2301 4317 2339 4323
rect 93 4297 131 4303
rect 429 4297 467 4303
rect 532 4297 563 4303
rect 621 4297 636 4303
rect 13 4277 51 4283
rect 221 4283 227 4296
rect 205 4277 227 4283
rect 205 4257 211 4277
rect 269 4277 323 4283
rect 621 4277 627 4297
rect 669 4297 723 4303
rect 1021 4297 1052 4303
rect 1085 4297 1100 4303
rect 1300 4297 1315 4303
rect 1373 4297 1404 4303
rect 1421 4297 1475 4303
rect 1645 4297 1708 4303
rect 1548 4292 1556 4296
rect 1828 4297 1843 4303
rect 1924 4297 1939 4303
rect 1949 4297 1964 4303
rect 2125 4297 2147 4303
rect 2564 4297 2595 4303
rect 2733 4303 2739 4323
rect 3405 4317 3420 4323
rect 2708 4297 2739 4303
rect 2749 4297 2780 4303
rect 2964 4297 2979 4303
rect 3028 4297 3043 4303
rect 3156 4297 3187 4303
rect 3789 4297 3804 4303
rect 3853 4303 3859 4323
rect 4893 4317 4915 4323
rect 3821 4297 3859 4303
rect 3869 4297 3907 4303
rect 3997 4297 4051 4303
rect 4061 4297 4076 4303
rect 4196 4297 4211 4303
rect 4573 4297 4588 4303
rect 4852 4297 4867 4303
rect 4877 4297 4892 4303
rect 5508 4297 5523 4303
rect 5741 4303 5747 4323
rect 5741 4297 5779 4303
rect 6045 4303 6051 4323
rect 6324 4316 6332 4324
rect 6388 4317 6419 4323
rect 6941 4317 6979 4323
rect 7284 4317 7299 4323
rect 7332 4316 7340 4324
rect 7396 4316 7404 4324
rect 7421 4317 7443 4323
rect 6013 4297 6051 4303
rect 6541 4297 6563 4303
rect 6828 4303 6836 4308
rect 6813 4297 6836 4303
rect 925 4277 940 4283
rect 1252 4277 1283 4283
rect 1309 4277 1347 4283
rect 2333 4277 2355 4283
rect 3773 4277 3788 4283
rect 4170 4276 4172 4284
rect 4525 4277 4547 4283
rect 4804 4277 4851 4283
rect 5677 4277 5699 4283
rect 5869 4277 5923 4283
rect 6813 4277 6819 4297
rect 7508 4297 7523 4303
rect 7796 4297 7811 4303
rect 8077 4297 8092 4303
rect 7192 4276 7196 4284
rect 7460 4277 7475 4283
rect 7485 4277 7539 4283
rect 7645 4277 7667 4283
rect 7725 4277 7763 4283
rect 8125 4277 8140 4283
rect 1868 4264 1876 4272
rect 2941 4257 2963 4263
rect 5940 4257 5955 4263
rect 6420 4256 6428 4264
rect 7996 4263 8004 4272
rect 7972 4257 8004 4263
rect 372 4236 374 4244
rect 1204 4236 1206 4244
rect 4388 4236 4392 4244
rect 5076 4236 5080 4244
rect 6852 4237 6867 4243
rect 8106 4236 8108 4244
rect 3272 4206 3278 4214
rect 3286 4206 3292 4214
rect 3300 4206 3306 4214
rect 3314 4206 3320 4214
rect 6344 4206 6350 4214
rect 6358 4206 6364 4214
rect 6372 4206 6378 4214
rect 6386 4206 6392 4214
rect 2104 4176 2108 4184
rect 2573 4177 2588 4183
rect 2872 4176 2876 4184
rect 6136 4176 6140 4184
rect 6442 4176 6444 4184
rect 7048 4176 7052 4184
rect 7226 4176 7228 4184
rect 7754 4176 7756 4184
rect 1229 4157 1252 4163
rect 1244 4154 1252 4157
rect 316 4143 324 4148
rect 860 4144 868 4148
rect 301 4137 324 4143
rect 1197 4137 1219 4143
rect 1540 4137 1555 4143
rect 1588 4137 1603 4143
rect 1636 4137 1667 4143
rect 1693 4137 1747 4143
rect 1837 4137 1868 4143
rect 2029 4143 2035 4163
rect 2477 4157 2492 4163
rect 2029 4137 2044 4143
rect 2196 4137 2211 4143
rect 589 4117 611 4123
rect 941 4117 979 4123
rect 973 4097 979 4117
rect 1181 4117 1196 4123
rect 1485 4117 1500 4123
rect 2317 4117 2332 4123
rect 2621 4123 2627 4143
rect 3037 4143 3043 4163
rect 4356 4157 4371 4163
rect 4813 4157 4860 4163
rect 5357 4157 5395 4163
rect 8084 4157 8115 4163
rect 2996 4137 3011 4143
rect 3037 4137 3052 4143
rect 3165 4137 3180 4143
rect 3220 4137 3235 4143
rect 3645 4137 3667 4143
rect 4268 4143 4276 4148
rect 4268 4137 4291 4143
rect 4301 4137 4316 4143
rect 4852 4137 4883 4143
rect 5405 4137 5443 4143
rect 2604 4117 2627 4123
rect 2604 4112 2612 4117
rect 3085 4117 3107 4123
rect 3213 4117 3251 4123
rect 3476 4117 3491 4123
rect 4013 4117 4051 4123
rect 989 4097 1004 4103
rect 1581 4097 1619 4103
rect 1940 4097 1955 4103
rect 1965 4097 1987 4103
rect 2173 4097 2188 4103
rect 3853 4097 3875 4103
rect 4045 4097 4051 4117
rect 4445 4117 4467 4123
rect 4500 4117 4531 4123
rect 4685 4117 4716 4123
rect 4724 4117 4755 4123
rect 4788 4117 4803 4123
rect 4941 4117 4995 4123
rect 5165 4117 5187 4123
rect 5437 4117 5443 4137
rect 5709 4137 5740 4143
rect 7149 4137 7180 4143
rect 7693 4137 7708 4143
rect 7780 4137 7788 4143
rect 8100 4137 8131 4143
rect 5501 4117 5516 4123
rect 5597 4117 5635 4123
rect 5789 4117 5811 4123
rect 5549 4097 5564 4103
rect 5597 4097 5603 4117
rect 6493 4117 6547 4123
rect 6573 4117 6611 4123
rect 6621 4117 6643 4123
rect 5677 4097 5692 4103
rect 6573 4097 6579 4117
rect 6900 4117 6915 4123
rect 7117 4117 7139 4123
rect 7293 4117 7324 4123
rect 7421 4117 7459 4123
rect 7501 4117 7523 4123
rect 7533 4117 7548 4123
rect 6756 4096 6764 4104
rect 7316 4097 7331 4103
rect 7421 4097 7427 4117
rect 7597 4117 7612 4123
rect 7796 4117 7811 4123
rect 7725 4097 7747 4103
rect 7908 4097 7923 4103
rect 3260 4083 3268 4088
rect 7740 4084 7748 4088
rect 8092 4084 8100 4088
rect 3260 4077 3308 4083
rect 4548 4077 4579 4083
rect 4573 4057 4579 4077
rect 6934 4076 6940 4084
rect 7885 4077 7900 4083
rect 7885 4057 7891 4077
rect 8020 4077 8035 4083
rect 36 4036 38 4044
rect 3828 4036 3830 4044
rect 4474 4036 4476 4044
rect 7354 4036 7356 4044
rect 7812 4036 7814 4044
rect 7946 4036 7948 4044
rect 1736 4006 1742 4014
rect 1750 4006 1756 4014
rect 1764 4006 1770 4014
rect 1778 4006 1784 4014
rect 4808 4006 4814 4014
rect 4822 4006 4828 4014
rect 4836 4006 4842 4014
rect 4850 4006 4856 4014
rect 740 3976 742 3984
rect 2388 3976 2390 3984
rect 3060 3976 3062 3984
rect 5226 3976 5228 3984
rect 8042 3976 8044 3984
rect 948 3956 952 3964
rect 6676 3936 6682 3944
rect 476 3932 484 3936
rect 2316 3932 2324 3936
rect 4892 3932 4900 3936
rect 269 3917 292 3923
rect 284 3912 292 3917
rect 765 3903 771 3923
rect 765 3897 803 3903
rect 1069 3903 1075 3923
rect 2740 3917 2771 3923
rect 3613 3917 3628 3923
rect 3748 3916 3756 3924
rect 4765 3917 4787 3923
rect 5309 3917 5324 3923
rect 5716 3916 5724 3924
rect 5828 3917 5843 3923
rect 6900 3916 6908 3924
rect 1037 3897 1075 3903
rect 1501 3897 1516 3903
rect 1636 3897 1651 3903
rect 1876 3897 1891 3903
rect 2493 3897 2508 3903
rect 2612 3897 2627 3903
rect 2765 3897 2787 3903
rect 3204 3897 3219 3903
rect 3485 3897 3500 3903
rect 3668 3897 3683 3903
rect 3693 3897 3724 3903
rect 5181 3897 5196 3903
rect 5501 3897 5532 3903
rect 5677 3897 5715 3903
rect 5748 3897 5779 3903
rect 6724 3897 6755 3903
rect 7364 3897 7395 3903
rect 8076 3903 8084 3908
rect 8061 3897 8084 3903
rect 1677 3877 1699 3883
rect 1828 3877 1843 3883
rect 1981 3877 2003 3883
rect 2237 3877 2259 3883
rect 2477 3877 2492 3883
rect 2692 3877 2723 3883
rect 2813 3877 2828 3883
rect 3357 3877 3411 3883
rect 3501 3877 3516 3883
rect 573 3857 595 3863
rect 1709 3857 1756 3863
rect 2204 3863 2212 3866
rect 2204 3857 2227 3863
rect 2580 3857 2595 3863
rect 3501 3857 3507 3877
rect 3645 3877 3667 3883
rect 4109 3877 4131 3883
rect 5245 3877 5283 3883
rect 6253 3877 6275 3883
rect 6557 3877 6579 3883
rect 6925 3877 6947 3883
rect 7357 3877 7372 3883
rect 8061 3877 8067 3897
rect 4884 3857 4915 3863
rect 5908 3856 5916 3864
rect 6972 3863 6980 3866
rect 6957 3857 6980 3863
rect 260 3836 262 3844
rect 490 3836 492 3844
rect 1732 3837 1779 3843
rect 4676 3837 4691 3843
rect 3272 3806 3278 3814
rect 3286 3806 3292 3814
rect 3300 3806 3306 3814
rect 3314 3806 3320 3814
rect 6344 3806 6350 3814
rect 6358 3806 6364 3814
rect 6372 3806 6378 3814
rect 6386 3806 6392 3814
rect 2532 3776 2534 3784
rect 2970 3776 2972 3784
rect 6013 3777 6028 3783
rect 6554 3776 6556 3784
rect 932 3756 940 3764
rect 1197 3757 1235 3763
rect 2132 3756 2140 3764
rect 2324 3756 2332 3764
rect 2637 3757 2659 3763
rect 4836 3757 4883 3763
rect 6132 3756 6140 3764
rect 221 3737 243 3743
rect 580 3737 611 3743
rect 708 3737 732 3743
rect 877 3737 931 3743
rect 1181 3737 1196 3743
rect 1453 3737 1484 3743
rect 2429 3737 2444 3743
rect 2637 3737 2652 3743
rect 3604 3737 3619 3743
rect 3693 3737 3708 3743
rect 3981 3737 4003 3743
rect 5005 3737 5043 3743
rect 5469 3737 5491 3743
rect 5773 3737 5788 3743
rect 5821 3737 5836 3743
rect 6500 3737 6531 3743
rect 6557 3737 6611 3743
rect 6733 3737 6748 3743
rect 6765 3743 6771 3763
rect 6973 3757 6996 3763
rect 6988 3754 6996 3757
rect 6765 3737 6780 3743
rect 6797 3737 6851 3743
rect 7389 3737 7411 3743
rect 7565 3737 7619 3743
rect 7709 3737 7731 3743
rect 7837 3737 7868 3743
rect 7924 3737 7940 3743
rect 77 3717 92 3723
rect 532 3717 563 3723
rect 852 3717 867 3723
rect 1149 3717 1171 3723
rect 1501 3717 1532 3723
rect 1581 3717 1596 3723
rect 156 3704 164 3714
rect 605 3697 627 3703
rect 1581 3697 1587 3717
rect 1661 3717 1699 3723
rect 2148 3717 2179 3723
rect 2189 3717 2220 3723
rect 2541 3717 2579 3723
rect 2141 3697 2147 3716
rect 2541 3697 2547 3717
rect 2669 3717 2684 3723
rect 2845 3717 2860 3723
rect 2845 3697 2851 3717
rect 3261 3717 3276 3723
rect 3965 3717 3980 3723
rect 4237 3717 4259 3723
rect 4380 3723 4388 3728
rect 4380 3717 4396 3723
rect 4628 3717 4643 3723
rect 4676 3717 4691 3723
rect 4797 3717 4828 3723
rect 4941 3717 4979 3723
rect 4973 3697 4979 3717
rect 6029 3704 6035 3723
rect 6164 3717 6195 3723
rect 6205 3717 6227 3723
rect 6333 3717 6419 3723
rect 5853 3697 5875 3703
rect 6349 3697 6396 3703
rect 6413 3697 6419 3717
rect 6717 3717 6732 3723
rect 7485 3717 7523 3723
rect 7661 3717 7692 3723
rect 7732 3717 7747 3723
rect 7773 3717 7811 3723
rect 7773 3697 7779 3717
rect 7844 3717 7859 3723
rect 477 3677 492 3683
rect 1052 3683 1060 3688
rect 1044 3677 1060 3683
rect 2316 3684 2324 3688
rect 3204 3677 3219 3683
rect 3596 3683 3604 3688
rect 6908 3684 6916 3688
rect 3596 3677 3612 3683
rect 6013 3677 6044 3683
rect 3258 3656 3260 3664
rect 820 3636 822 3644
rect 3434 3636 3436 3644
rect 5962 3636 5964 3644
rect 6084 3636 6086 3644
rect 1736 3606 1742 3614
rect 1750 3606 1756 3614
rect 1764 3606 1770 3614
rect 1778 3606 1784 3614
rect 4808 3606 4814 3614
rect 4822 3606 4828 3614
rect 4836 3606 4842 3614
rect 4850 3606 4856 3614
rect 1098 3556 1100 3564
rect 3802 3556 3804 3564
rect 7002 3556 7004 3564
rect 2660 3537 2691 3543
rect 5732 3536 5734 3544
rect 5908 3537 5923 3543
rect 6388 3537 6435 3543
rect 6508 3537 6524 3543
rect 5084 3532 5092 3536
rect 205 3497 227 3503
rect 285 3497 307 3503
rect 413 3497 435 3503
rect 1069 3503 1075 3523
rect 2276 3516 2284 3524
rect 1133 3503 1139 3516
rect 1012 3497 1027 3503
rect 1037 3497 1075 3503
rect 1101 3497 1139 3503
rect 1149 3497 1203 3503
rect 1236 3497 1251 3503
rect 1684 3497 1715 3503
rect 2365 3503 2371 3523
rect 3293 3517 3356 3523
rect 3373 3517 3388 3523
rect 3549 3517 3587 3523
rect 3725 3517 3763 3523
rect 2333 3497 2371 3503
rect 2381 3497 2419 3503
rect 2525 3497 2540 3503
rect 2829 3497 2851 3503
rect 3709 3497 3740 3503
rect 3757 3497 3772 3503
rect 4004 3497 4019 3503
rect 4372 3497 4403 3503
rect 4413 3497 4467 3503
rect 4564 3497 4579 3503
rect 4589 3497 4604 3503
rect 4733 3503 4739 3523
rect 5012 3517 5027 3523
rect 5549 3517 5571 3523
rect 5620 3516 5628 3524
rect 4685 3497 4723 3503
rect 4733 3497 4771 3503
rect 5165 3497 5196 3503
rect 5508 3497 5523 3503
rect 5533 3497 5548 3503
rect 5652 3497 5683 3503
rect 5700 3497 5731 3503
rect 5869 3497 5891 3503
rect 6724 3497 6739 3503
rect 6973 3503 6979 3523
rect 6941 3497 6979 3503
rect 7005 3497 7020 3503
rect 7037 3503 7043 3523
rect 7133 3517 7148 3523
rect 7028 3497 7043 3503
rect 7053 3497 7107 3503
rect 7229 3497 7251 3503
rect 7741 3503 7747 3523
rect 7709 3497 7747 3503
rect 349 3477 387 3483
rect 381 3457 387 3477
rect 1380 3476 1384 3484
rect 1485 3477 1539 3483
rect 1773 3477 1788 3483
rect 2237 3477 2259 3483
rect 2461 3477 2515 3483
rect 2612 3477 2643 3483
rect 2653 3477 2675 3483
rect 2685 3477 2707 3483
rect 2060 3463 2068 3472
rect 2669 3464 2675 3477
rect 3405 3477 3459 3483
rect 3624 3476 3628 3484
rect 3852 3477 3868 3483
rect 3852 3476 3860 3477
rect 4349 3477 4364 3483
rect 4605 3477 4620 3483
rect 4781 3477 4796 3483
rect 4941 3477 4995 3483
rect 5044 3477 5059 3483
rect 5565 3477 5603 3483
rect 5700 3477 5715 3483
rect 6429 3477 6467 3483
rect 6541 3477 6563 3483
rect 6860 3477 6876 3483
rect 6860 3476 6868 3477
rect 2060 3457 2092 3463
rect 4317 3457 4332 3463
rect 6077 3457 6092 3463
rect 6340 3456 6348 3464
rect 1482 3436 1484 3444
rect 3293 3437 3340 3443
rect 3540 3436 3542 3444
rect 5076 3436 5078 3444
rect 5386 3436 5388 3444
rect 6154 3436 6156 3444
rect 7754 3436 7756 3444
rect 3272 3406 3278 3414
rect 3286 3406 3292 3414
rect 3300 3406 3306 3414
rect 3314 3406 3320 3414
rect 6344 3406 6350 3414
rect 6358 3406 6364 3414
rect 6372 3406 6378 3414
rect 6386 3406 6392 3414
rect 100 3377 115 3383
rect 3293 3377 3340 3383
rect 4680 3376 4684 3384
rect 4836 3377 4883 3383
rect 5428 3376 5430 3384
rect 6522 3376 6524 3384
rect 6596 3376 6600 3384
rect 6968 3376 6972 3384
rect 173 3337 188 3343
rect 365 3343 371 3363
rect 356 3337 371 3343
rect 877 3343 883 3363
rect 6404 3357 6419 3363
rect 845 3337 867 3343
rect 877 3337 892 3343
rect 909 3337 963 3343
rect 1012 3337 1027 3343
rect 1764 3337 1827 3343
rect 1901 3337 1923 3343
rect 2804 3337 2819 3343
rect 2893 3337 2915 3343
rect 3348 3337 3363 3343
rect 3437 3337 3459 3343
rect 3821 3337 3852 3343
rect 3892 3337 3907 3343
rect 4941 3343 4947 3356
rect 4925 3337 4947 3343
rect 5245 3337 5283 3343
rect 5469 3337 5500 3343
rect 5661 3343 5667 3356
rect 5645 3337 5667 3343
rect 5677 3337 5699 3343
rect 6172 3343 6180 3348
rect 6116 3337 6147 3343
rect 6157 3337 6180 3343
rect 7005 3337 7020 3343
rect 7597 3343 7603 3356
rect 7597 3337 7619 3343
rect 8141 3337 8156 3343
rect 381 3317 396 3323
rect 621 3317 659 3323
rect 621 3297 627 3317
rect 861 3317 892 3323
rect 1053 3317 1068 3323
rect 1341 3317 1363 3323
rect 1885 3317 1900 3323
rect 3244 3324 3252 3328
rect 2525 3317 2540 3323
rect 2669 3317 2723 3323
rect 2765 3317 2803 3323
rect 3869 3317 3891 3323
rect 3924 3317 3955 3323
rect 5300 3317 5315 3323
rect 5373 3317 5404 3323
rect 5629 3317 5660 3323
rect 5725 3317 5763 3323
rect 2605 3297 2643 3303
rect 2868 3296 2876 3304
rect 4068 3296 4072 3304
rect 84 3277 115 3283
rect 292 3276 296 3284
rect 2134 3276 2140 3284
rect 3405 3277 3420 3283
rect 3693 3277 3708 3283
rect 5021 3283 5027 3303
rect 5277 3297 5299 3303
rect 5757 3297 5763 3317
rect 6093 3317 6131 3323
rect 6716 3324 6724 3328
rect 6461 3317 6483 3323
rect 6125 3297 6131 3317
rect 7101 3317 7123 3323
rect 7229 3317 7251 3323
rect 7773 3317 7827 3323
rect 8013 3317 8035 3323
rect 6372 3297 6419 3303
rect 7581 3297 7596 3303
rect 7764 3296 7772 3304
rect 5005 3277 5027 3283
rect 5226 3276 5228 3284
rect 7700 3276 7702 3284
rect 5786 3256 5788 3264
rect 826 3236 828 3244
rect 2724 3236 2726 3244
rect 5108 3236 5110 3244
rect 1736 3206 1742 3214
rect 1750 3206 1756 3214
rect 1764 3206 1770 3214
rect 1778 3206 1784 3214
rect 4808 3206 4814 3214
rect 4822 3206 4828 3214
rect 4836 3206 4842 3214
rect 4850 3206 4856 3214
rect 740 3176 742 3184
rect 1482 3176 1484 3184
rect 4564 3176 4566 3184
rect 4900 3176 4902 3184
rect 5050 3176 5052 3184
rect 6986 3156 6988 3164
rect 44 3137 60 3143
rect 44 3132 52 3137
rect 3460 3136 3462 3144
rect 3924 3136 3930 3144
rect 1228 3132 1236 3136
rect 2012 3132 2020 3136
rect 5772 3132 5780 3136
rect 488 3116 492 3124
rect 1380 3117 1411 3123
rect 1421 3117 1459 3123
rect 1597 3117 1612 3123
rect 372 3097 387 3103
rect 589 3097 611 3103
rect 820 3097 835 3103
rect 1117 3097 1148 3103
rect 1309 3097 1363 3103
rect 1485 3097 1532 3103
rect 1725 3097 1740 3103
rect 1869 3103 1875 3123
rect 2372 3116 2380 3124
rect 1764 3097 1795 3103
rect 1869 3097 1907 3103
rect 2061 3097 2099 3103
rect 2397 3103 2403 3123
rect 2836 3116 2840 3124
rect 3181 3117 3196 3123
rect 2397 3097 2435 3103
rect 3309 3097 3324 3103
rect 3485 3103 3491 3123
rect 3485 3097 3523 3103
rect 3629 3097 3644 3103
rect 3725 3103 3731 3123
rect 3837 3117 3852 3123
rect 3684 3097 3715 3103
rect 3725 3097 3763 3103
rect 3988 3097 4003 3103
rect 4285 3097 4300 3103
rect 4589 3103 4595 3123
rect 4589 3097 4627 3103
rect 4685 3097 4739 3103
rect 5021 3097 5043 3103
rect 5373 3097 5395 3103
rect 5453 3097 5475 3103
rect 6180 3097 6195 3103
rect 6333 3103 6339 3123
rect 6333 3097 6419 3103
rect 6621 3097 6668 3103
rect 6876 3103 6884 3108
rect 6876 3097 6899 3103
rect 29 3077 60 3083
rect 269 3077 284 3083
rect 269 3057 275 3077
rect 797 3077 851 3083
rect 1325 3077 1340 3083
rect 1629 3077 1683 3083
rect 2020 3077 2051 3083
rect 2333 3077 2355 3083
rect 2541 3077 2572 3083
rect 3572 3077 3587 3083
rect 3636 3077 3667 3083
rect 3844 3077 3875 3083
rect 5100 3077 5116 3083
rect 5100 3076 5108 3077
rect 5549 3077 5564 3083
rect 6516 3077 6531 3083
rect 6557 3077 6611 3083
rect 6893 3077 6899 3097
rect 6957 3103 6963 3123
rect 7069 3117 7084 3123
rect 7108 3116 7116 3124
rect 7908 3116 7916 3124
rect 6925 3097 6963 3103
rect 7117 3097 7171 3103
rect 7188 3097 7203 3103
rect 8036 3097 8067 3103
rect 7677 3077 7699 3083
rect 2004 3057 2035 3063
rect 2660 3056 2668 3064
rect 4797 3057 4883 3063
rect 7037 3057 7052 3063
rect 7228 3063 7236 3066
rect 7677 3064 7683 3077
rect 8026 3076 8028 3084
rect 7213 3057 7236 3063
rect 7444 3056 7452 3064
rect 116 3036 118 3044
rect 1242 3036 1244 3044
rect 2596 3036 2598 3044
rect 6554 3036 6556 3044
rect 6772 3036 6774 3044
rect 7716 3036 7718 3044
rect 3272 3006 3278 3014
rect 3286 3006 3292 3014
rect 3300 3006 3306 3014
rect 3314 3006 3320 3014
rect 6344 3006 6350 3014
rect 6358 3006 6364 3014
rect 6372 3006 6378 3014
rect 6386 3006 6392 3014
rect 2372 2976 2374 2984
rect 3309 2977 3331 2983
rect 1324 2957 1347 2963
rect 1324 2954 1332 2957
rect 2228 2957 2260 2963
rect 2252 2948 2260 2957
rect 3309 2963 3315 2977
rect 3482 2976 3484 2984
rect 3720 2976 3724 2984
rect 6285 2977 6316 2983
rect 3261 2957 3315 2963
rect 5181 2957 5228 2963
rect 5565 2957 5587 2963
rect 52 2937 67 2943
rect 109 2937 131 2943
rect 260 2937 275 2943
rect 1677 2937 1699 2943
rect 1812 2937 1843 2943
rect 1869 2937 1884 2943
rect 1949 2937 1971 2943
rect 2061 2937 2083 2943
rect 2477 2937 2531 2943
rect 2580 2937 2595 2943
rect 2957 2937 2979 2943
rect 3245 2937 3324 2943
rect 3869 2937 3907 2943
rect 237 2917 259 2923
rect 317 2917 355 2923
rect 445 2917 460 2923
rect 212 2896 220 2904
rect 237 2897 243 2917
rect 829 2917 867 2923
rect 829 2897 835 2917
rect 1597 2917 1635 2923
rect 1629 2897 1635 2917
rect 1812 2917 1827 2923
rect 1997 2917 2012 2923
rect 2637 2917 2675 2923
rect 2669 2897 2675 2917
rect 3213 2917 3235 2923
rect 3389 2917 3427 2923
rect 3789 2917 3820 2923
rect 4029 2917 4067 2923
rect 4004 2896 4012 2904
rect 4029 2897 4035 2917
rect 4093 2923 4099 2943
rect 4669 2937 4723 2943
rect 4781 2937 4819 2943
rect 4093 2917 4116 2923
rect 4108 2912 4116 2917
rect 4461 2917 4499 2923
rect 4461 2897 4467 2917
rect 4813 2923 4819 2937
rect 5261 2943 5267 2956
rect 7548 2944 7556 2948
rect 5245 2937 5267 2943
rect 5692 2943 5700 2944
rect 5629 2937 5651 2943
rect 5692 2937 5708 2943
rect 5784 2936 5788 2944
rect 7044 2937 7059 2943
rect 7805 2937 7827 2943
rect 4813 2917 4904 2923
rect 5908 2917 5923 2923
rect 6100 2917 6115 2923
rect 6557 2917 6572 2923
rect 6877 2917 6915 2923
rect 6877 2897 6883 2917
rect 7021 2917 7036 2923
rect 7140 2917 7171 2923
rect 7421 2917 7452 2923
rect 7421 2897 7427 2917
rect 7636 2917 7651 2923
rect 7844 2896 7852 2904
rect 5212 2884 5220 2888
rect 1286 2876 1292 2884
rect 1956 2877 1971 2883
rect 4358 2876 4364 2884
rect 5028 2877 5043 2883
rect 5748 2877 5779 2883
rect 6676 2876 6682 2884
rect 7524 2877 7539 2883
rect 8109 2877 8156 2883
rect 1736 2806 1742 2814
rect 1750 2806 1756 2814
rect 1764 2806 1770 2814
rect 1778 2806 1784 2814
rect 4808 2806 4814 2814
rect 4822 2806 4828 2814
rect 4836 2806 4842 2814
rect 4850 2806 4856 2814
rect 3252 2777 3267 2783
rect 5828 2776 5830 2784
rect 4762 2756 4764 2764
rect 748 2732 756 2736
rect 1382 2736 1388 2744
rect 5524 2737 5539 2743
rect 5690 2736 5692 2744
rect 6212 2736 6218 2744
rect 7789 2737 7812 2743
rect 7972 2736 7974 2744
rect 8077 2737 8092 2743
rect 892 2732 900 2736
rect 4796 2732 4804 2736
rect 420 2716 428 2724
rect 1172 2716 1176 2724
rect 1604 2716 1612 2724
rect 1780 2717 1795 2723
rect 1965 2717 1987 2723
rect 900 2697 915 2703
rect 973 2697 995 2703
rect 1636 2697 1667 2703
rect 1677 2697 1692 2703
rect 1828 2697 1859 2703
rect 2180 2696 2184 2704
rect 3501 2697 3523 2703
rect 3588 2697 3640 2703
rect 3821 2703 3827 2723
rect 3773 2697 3811 2703
rect 3821 2697 3859 2703
rect 3949 2697 3964 2703
rect 4333 2703 4339 2723
rect 5421 2717 5459 2723
rect 4301 2697 4339 2703
rect 4349 2697 4387 2703
rect 4564 2697 4579 2703
rect 5373 2697 5411 2703
rect 5661 2703 5667 2723
rect 5604 2697 5619 2703
rect 5629 2697 5667 2703
rect 5757 2697 5772 2703
rect 6093 2703 6099 2723
rect 6052 2697 6067 2703
rect 6093 2697 6131 2703
rect 6276 2697 6291 2703
rect 7229 2703 7235 2723
rect 7197 2697 7235 2703
rect 7812 2697 7827 2703
rect 445 2677 467 2683
rect 484 2677 499 2683
rect 1693 2677 1715 2683
rect 1821 2677 1836 2683
rect 1933 2677 1948 2683
rect 3133 2677 3155 2683
rect 3508 2677 3523 2683
rect 3581 2677 3596 2683
rect 4388 2677 4403 2683
rect 4429 2677 4483 2683
rect 4525 2677 4556 2683
rect 5101 2677 5123 2683
rect 5188 2677 5203 2683
rect 5277 2677 5331 2683
rect 5789 2677 5811 2683
rect 6029 2677 6051 2683
rect 7066 2676 7068 2684
rect 7277 2677 7299 2683
rect 7492 2677 7507 2683
rect 1404 2672 1412 2676
rect 1796 2656 1804 2664
rect 1949 2657 1955 2676
rect 1988 2656 1996 2664
rect 4781 2657 4812 2663
rect 5764 2657 5779 2663
rect 1108 2636 1110 2644
rect 3562 2636 3564 2644
rect 6452 2636 6456 2644
rect 3272 2606 3278 2614
rect 3286 2606 3292 2614
rect 3300 2606 3306 2614
rect 3314 2606 3320 2614
rect 6344 2606 6350 2614
rect 6358 2606 6364 2614
rect 6372 2606 6378 2614
rect 6386 2606 6392 2614
rect 5236 2576 5238 2584
rect 6052 2576 6054 2584
rect 1213 2557 1228 2563
rect 2237 2557 2275 2563
rect 3932 2557 3964 2563
rect 3932 2548 3940 2557
rect 765 2537 796 2543
rect 1108 2537 1123 2543
rect 1293 2537 1308 2543
rect 1373 2537 1427 2543
rect 2429 2537 2451 2543
rect 3316 2537 3379 2543
rect 4301 2543 4307 2556
rect 4237 2537 4291 2543
rect 4301 2537 4323 2543
rect 5197 2543 5203 2563
rect 5197 2537 5212 2543
rect 5373 2537 5395 2543
rect 5837 2543 5843 2563
rect 6301 2557 6323 2563
rect 7661 2557 7676 2563
rect 5789 2537 5827 2543
rect 5837 2537 5852 2543
rect 6717 2537 6739 2543
rect 7245 2537 7267 2543
rect 7677 2537 7699 2543
rect 852 2517 883 2523
rect 900 2517 915 2523
rect 973 2517 1027 2523
rect 1245 2517 1260 2523
rect 1988 2517 2019 2523
rect 2029 2517 2051 2523
rect 2301 2517 2323 2523
rect 2413 2517 2428 2523
rect 2605 2517 2627 2523
rect 2877 2517 2931 2523
rect 3021 2517 3059 2523
rect 3069 2517 3123 2523
rect 932 2497 947 2503
rect 964 2496 972 2504
rect 1277 2497 1315 2503
rect 1325 2497 1340 2503
rect 1981 2497 1987 2516
rect 2372 2497 2387 2503
rect 3021 2497 3027 2517
rect 3517 2517 3555 2523
rect 3405 2497 3420 2503
rect 3549 2497 3555 2517
rect 3716 2517 3731 2523
rect 4333 2517 4371 2523
rect 4365 2497 4371 2517
rect 5044 2517 5059 2523
rect 5245 2517 5276 2523
rect 5165 2497 5187 2503
rect 5245 2497 5251 2517
rect 5293 2517 5331 2523
rect 5325 2497 5331 2517
rect 5460 2517 5475 2523
rect 5597 2517 5635 2523
rect 5677 2517 5692 2523
rect 5549 2497 5564 2503
rect 5597 2497 5603 2517
rect 5821 2517 5852 2523
rect 5997 2517 6028 2523
rect 6221 2517 6252 2523
rect 6308 2517 6323 2523
rect 7165 2517 7203 2523
rect 6189 2497 6204 2503
rect 7197 2497 7203 2517
rect 7229 2517 7244 2523
rect 7677 2524 7683 2537
rect 7748 2517 7779 2523
rect 7853 2517 7875 2523
rect 7997 2517 8012 2523
rect 8036 2517 8051 2523
rect 7773 2497 7804 2503
rect 4620 2484 4628 2488
rect 3578 2476 3580 2484
rect 4404 2477 4419 2483
rect 4532 2477 4556 2483
rect 5412 2477 5427 2483
rect 1658 2456 1660 2464
rect 1066 2436 1068 2444
rect 2292 2436 2294 2444
rect 2634 2436 2636 2444
rect 6106 2436 6108 2444
rect 1736 2406 1742 2414
rect 1750 2406 1756 2414
rect 1764 2406 1770 2414
rect 1778 2406 1784 2414
rect 4808 2406 4814 2414
rect 4822 2406 4828 2414
rect 4836 2406 4842 2414
rect 4850 2406 4856 2414
rect 7476 2376 7478 2384
rect 516 2356 518 2364
rect 7338 2356 7340 2364
rect 2842 2336 2844 2344
rect 5837 2337 5875 2343
rect 1516 2332 1524 2336
rect 4508 2332 4516 2336
rect 548 2297 579 2303
rect 589 2297 604 2303
rect 717 2297 732 2303
rect 1421 2297 1459 2303
rect 1908 2297 1923 2303
rect 2068 2297 2083 2303
rect 2349 2297 2371 2303
rect 2701 2297 2716 2303
rect 2813 2303 2819 2323
rect 2932 2317 2947 2323
rect 4493 2317 4515 2323
rect 2781 2297 2819 2303
rect 2973 2297 3027 2303
rect 3181 2297 3203 2303
rect 3213 2297 3228 2303
rect 3293 2297 3340 2303
rect 4717 2303 4723 2323
rect 4852 2317 4899 2323
rect 4685 2297 4723 2303
rect 5092 2297 5144 2303
rect 5421 2297 5475 2303
rect 5837 2297 5843 2337
rect 5924 2336 5926 2344
rect 5949 2317 5987 2323
rect 6045 2317 6060 2323
rect 5869 2297 5923 2303
rect 6132 2297 6147 2303
rect 6221 2297 6243 2303
rect 6349 2297 6419 2303
rect 6596 2297 6611 2303
rect 6957 2303 6963 2323
rect 6980 2316 6988 2324
rect 7572 2317 7596 2323
rect 6925 2297 6963 2303
rect 7309 2297 7331 2303
rect 7380 2297 7395 2303
rect 7508 2297 7539 2303
rect 7709 2303 7715 2323
rect 7677 2297 7715 2303
rect 8036 2297 8051 2303
rect 461 2277 499 2283
rect 1325 2277 1379 2283
rect 1476 2277 1491 2283
rect 1581 2277 1603 2283
rect 1997 2277 2019 2283
rect 3348 2277 3364 2283
rect 4029 2277 4051 2283
rect 5085 2277 5107 2283
rect 5197 2277 5219 2283
rect 5085 2264 5091 2277
rect 5981 2277 6003 2283
rect 6845 2277 6860 2283
rect 7005 2277 7027 2283
rect 7364 2277 7379 2283
rect 7437 2277 7452 2283
rect 1828 2257 1891 2263
rect 3229 2257 3251 2263
rect 5028 2256 5036 2264
rect 7373 2257 7379 2277
rect 7629 2277 7644 2283
rect 260 2236 262 2244
rect 436 2236 438 2244
rect 1508 2236 1510 2244
rect 1805 2237 1852 2243
rect 4522 2236 4524 2244
rect 4580 2237 4595 2243
rect 5700 2236 5702 2244
rect 6084 2237 6099 2243
rect 6788 2236 6790 2244
rect 6826 2236 6828 2244
rect 7258 2236 7260 2244
rect 7796 2237 7811 2243
rect 3272 2206 3278 2214
rect 3286 2206 3292 2214
rect 3300 2206 3306 2214
rect 3314 2206 3320 2214
rect 6344 2206 6350 2214
rect 6358 2206 6364 2214
rect 6372 2206 6378 2214
rect 6386 2206 6392 2214
rect 1380 2176 1382 2184
rect 2580 2176 2582 2184
rect 2932 2177 2947 2183
rect 3498 2176 3500 2184
rect 4010 2176 4012 2184
rect 4804 2177 4835 2183
rect 5626 2176 5628 2184
rect 5892 2176 5894 2184
rect 6168 2176 6172 2184
rect 6612 2176 6614 2184
rect 1485 2157 1500 2163
rect 205 2137 227 2143
rect 397 2137 412 2143
rect 484 2137 499 2143
rect 532 2137 547 2143
rect 596 2137 611 2143
rect 717 2143 723 2156
rect 701 2137 723 2143
rect 1245 2137 1267 2143
rect 1693 2143 1699 2163
rect 1869 2157 1907 2163
rect 1980 2148 1988 2156
rect 1396 2137 1411 2143
rect 1421 2137 1491 2143
rect 1677 2137 1699 2143
rect 1773 2137 1788 2143
rect 77 2117 108 2123
rect 333 2117 371 2123
rect 381 2117 396 2123
rect 333 2097 339 2117
rect 404 2117 419 2123
rect 477 2117 492 2123
rect 557 2117 595 2123
rect 676 2117 691 2123
rect 1676 2124 1684 2128
rect 1229 2117 1244 2123
rect 1613 2117 1635 2123
rect 1773 2123 1779 2137
rect 3028 2137 3043 2143
rect 3917 2137 3939 2143
rect 4764 2137 4780 2143
rect 5501 2137 5555 2143
rect 5677 2143 5683 2163
rect 5677 2137 5692 2143
rect 6349 2137 6412 2143
rect 1725 2117 1779 2123
rect 1837 2117 1852 2123
rect 2164 2117 2195 2123
rect 3592 2116 3596 2124
rect 3725 2117 3747 2123
rect 3757 2117 3795 2123
rect 3821 2117 3875 2123
rect 3917 2117 3932 2123
rect 1389 2097 1404 2103
rect 2900 2097 2915 2103
rect 3789 2097 3795 2117
rect 4653 2117 4668 2123
rect 5229 2117 5260 2123
rect 5421 2117 5459 2123
rect 6493 2123 6499 2143
rect 6557 2137 6611 2143
rect 7101 2137 7116 2143
rect 7357 2137 7372 2143
rect 6476 2117 6499 2123
rect 6476 2112 6484 2117
rect 6701 2117 6739 2123
rect 3885 2097 3923 2103
rect 5373 2097 5411 2103
rect 5597 2097 5619 2103
rect 6733 2097 6739 2117
rect 6772 2117 6796 2123
rect 6941 2117 6963 2123
rect 7197 2117 7212 2123
rect 7373 2117 7396 2123
rect 7388 2114 7396 2117
rect 7844 2096 7852 2104
rect 3484 2084 3492 2088
rect 902 2076 908 2084
rect 1988 2076 1994 2084
rect 2724 2076 2726 2084
rect 3380 2077 3459 2083
rect 4068 2077 4083 2083
rect 6762 2076 6764 2084
rect 7789 2077 7804 2083
rect 8109 2077 8156 2083
rect 1604 2036 1606 2044
rect 1736 2006 1742 2014
rect 1750 2006 1756 2014
rect 1764 2006 1770 2014
rect 1778 2006 1784 2014
rect 4808 2006 4814 2014
rect 4822 2006 4828 2014
rect 4836 2006 4842 2014
rect 4850 2006 4856 2014
rect 3370 1976 3372 1984
rect 5178 1976 5180 1984
rect 3956 1956 3958 1964
rect 189 1937 204 1943
rect 724 1936 726 1944
rect 1242 1936 1244 1944
rect 2968 1936 2972 1944
rect 4712 1936 4716 1944
rect 5037 1937 5052 1943
rect 8109 1937 8156 1943
rect 276 1897 291 1903
rect 301 1897 323 1903
rect 204 1892 212 1896
rect 749 1903 755 1923
rect 916 1917 931 1923
rect 2253 1917 2268 1923
rect 708 1897 723 1903
rect 749 1897 787 1903
rect 1709 1897 1740 1903
rect 1988 1897 2003 1903
rect 2109 1897 2124 1903
rect 2365 1903 2371 1923
rect 2404 1916 2412 1924
rect 2301 1897 2355 1903
rect 2365 1897 2396 1903
rect 2429 1903 2435 1923
rect 2685 1917 2723 1923
rect 2756 1917 2771 1923
rect 3140 1916 3148 1924
rect 3252 1916 3260 1924
rect 3844 1917 3859 1923
rect 2429 1897 2467 1903
rect 2477 1897 2515 1903
rect 2532 1897 2547 1903
rect 3485 1897 3507 1903
rect 3981 1903 3987 1923
rect 3940 1897 3955 1903
rect 3981 1897 4019 1903
rect 4349 1903 4355 1923
rect 5108 1916 5116 1924
rect 5309 1917 5331 1923
rect 5684 1916 5692 1924
rect 4301 1897 4339 1903
rect 4349 1897 4387 1903
rect 4781 1897 4803 1903
rect 4813 1897 4860 1903
rect 5181 1897 5219 1903
rect 5325 1897 5379 1903
rect 5437 1897 5468 1903
rect 6349 1903 6355 1923
rect 7724 1917 7747 1923
rect 7724 1912 7732 1917
rect 7876 1916 7884 1924
rect 6349 1897 6435 1903
rect 6445 1897 6460 1903
rect 6500 1897 6515 1903
rect 6573 1897 6588 1903
rect 6621 1897 6643 1903
rect 7748 1897 7763 1903
rect 7901 1903 7907 1923
rect 7860 1897 7875 1903
rect 7901 1897 7916 1903
rect 8020 1897 8035 1903
rect 397 1877 419 1883
rect 973 1877 1027 1883
rect 1053 1877 1068 1883
rect 1101 1877 1155 1883
rect 1261 1877 1283 1883
rect 3101 1877 3123 1883
rect 3820 1877 3836 1883
rect 3820 1876 3828 1877
rect 4045 1877 4060 1883
rect 4077 1877 4131 1883
rect 4205 1877 4259 1883
rect 4749 1877 4764 1883
rect 4884 1877 4915 1883
rect 5517 1877 5539 1883
rect 6092 1877 6116 1883
rect 6212 1876 6214 1884
rect 6461 1877 6483 1883
rect 6580 1877 6611 1883
rect 6797 1877 6835 1883
rect 7373 1877 7395 1883
rect 7789 1877 7804 1883
rect 156 1864 164 1872
rect 3724 1863 3732 1866
rect 3724 1857 3747 1863
rect 4941 1857 4963 1863
rect 6628 1857 6643 1863
rect 2730 1836 2732 1844
rect 2778 1836 2780 1844
rect 3912 1836 3916 1844
rect 5300 1836 5302 1844
rect 6532 1836 6534 1844
rect 7818 1836 7820 1844
rect 7978 1836 7980 1844
rect 3272 1806 3278 1814
rect 3286 1806 3292 1814
rect 3300 1806 3306 1814
rect 3314 1806 3320 1814
rect 6344 1806 6350 1814
rect 6358 1806 6364 1814
rect 6372 1806 6378 1814
rect 6386 1806 6392 1814
rect 1034 1776 1036 1784
rect 2500 1776 2504 1784
rect 2788 1776 2790 1784
rect 6692 1776 6694 1784
rect 1773 1757 1827 1763
rect 493 1737 515 1743
rect 941 1737 956 1743
rect 1773 1743 1779 1757
rect 1972 1757 2004 1763
rect 1996 1748 2004 1757
rect 4980 1756 4988 1764
rect 6029 1757 6051 1763
rect 1757 1737 1779 1743
rect 2100 1737 2115 1743
rect 2125 1737 2163 1743
rect 2861 1737 2915 1743
rect 3085 1737 3139 1743
rect 3332 1737 3347 1743
rect 3412 1737 3427 1743
rect 3588 1737 3619 1743
rect 3661 1737 3699 1743
rect 3748 1737 3763 1743
rect 3860 1737 3875 1743
rect 4333 1737 4355 1743
rect 4916 1737 4963 1743
rect 5156 1737 5187 1743
rect 5532 1743 5540 1748
rect 5532 1737 5555 1743
rect 5565 1737 5596 1743
rect 5693 1737 5747 1743
rect 6909 1737 6931 1743
rect 7756 1737 7780 1743
rect 180 1717 195 1723
rect 205 1717 227 1723
rect 317 1717 332 1723
rect 452 1717 467 1723
rect 557 1717 579 1723
rect 589 1717 627 1723
rect 653 1717 707 1723
rect 125 1697 147 1703
rect 621 1697 627 1717
rect 804 1717 835 1723
rect 989 1717 1027 1723
rect 1021 1697 1027 1717
rect 1101 1717 1116 1723
rect 1332 1717 1347 1723
rect 1357 1717 1411 1723
rect 1741 1717 1804 1723
rect 2077 1717 2092 1723
rect 2973 1717 3011 1723
rect 2068 1696 2076 1704
rect 2724 1696 2732 1704
rect 3005 1697 3011 1717
rect 3389 1717 3404 1723
rect 3220 1697 3235 1703
rect 3389 1697 3395 1717
rect 3444 1717 3475 1723
rect 3485 1717 3500 1723
rect 3741 1717 3756 1723
rect 3885 1717 3923 1723
rect 3764 1697 3779 1703
rect 3828 1697 3843 1703
rect 3917 1697 3923 1717
rect 5021 1717 5107 1723
rect 5581 1717 5619 1723
rect 5581 1697 5587 1717
rect 5636 1717 5651 1723
rect 5997 1717 6019 1723
rect 6084 1717 6099 1723
rect 6244 1717 6259 1723
rect 6468 1717 6483 1723
rect 6765 1717 6803 1723
rect 6429 1697 6467 1703
rect 6701 1697 6723 1703
rect 6797 1697 6803 1717
rect 6932 1717 6947 1723
rect 6957 1717 6972 1723
rect 7092 1717 7107 1723
rect 7293 1717 7331 1723
rect 7325 1697 7331 1717
rect 141 1677 156 1683
rect 1116 1677 1139 1683
rect 1172 1676 1178 1684
rect 2140 1683 2148 1688
rect 4988 1684 4996 1688
rect 2029 1677 2052 1683
rect 2140 1677 2156 1683
rect 4442 1676 4444 1684
rect 4756 1676 4762 1684
rect 5036 1684 5044 1688
rect 6700 1684 6708 1688
rect 7212 1684 7220 1688
rect 7620 1676 7626 1684
rect 1684 1636 1686 1644
rect 3364 1636 3366 1644
rect 5988 1636 5990 1644
rect 6388 1637 6435 1643
rect 1736 1606 1742 1614
rect 1750 1606 1756 1614
rect 1764 1606 1770 1614
rect 1778 1606 1784 1614
rect 4808 1606 4814 1614
rect 4822 1606 4828 1614
rect 4836 1606 4842 1614
rect 4850 1606 4856 1614
rect 1956 1556 1960 1564
rect 52 1537 99 1543
rect 1236 1537 1252 1543
rect 1325 1537 1340 1543
rect 2541 1537 2564 1543
rect 2556 1532 2564 1537
rect 3596 1532 3604 1536
rect 4006 1536 4012 1544
rect 4212 1536 4214 1544
rect 6132 1536 6134 1544
rect 6845 1537 6860 1543
rect 7780 1536 7782 1544
rect 7908 1536 7910 1544
rect 3740 1532 3748 1536
rect 61 1517 76 1523
rect 205 1497 259 1503
rect 324 1497 339 1503
rect 461 1503 467 1523
rect 1172 1516 1180 1524
rect 2205 1517 2243 1523
rect 461 1497 483 1503
rect 580 1497 595 1503
rect 1156 1497 1171 1503
rect 1236 1497 1267 1503
rect 1277 1497 1331 1503
rect 2157 1497 2172 1503
rect 3821 1497 3843 1503
rect 4044 1503 4052 1506
rect 4044 1497 4067 1503
rect 4125 1497 4163 1503
rect 4237 1503 4243 1523
rect 5236 1516 5244 1524
rect 5677 1517 5692 1523
rect 5757 1517 5795 1523
rect 5812 1516 5820 1524
rect 6292 1517 6307 1523
rect 6404 1517 6419 1523
rect 6797 1517 6835 1523
rect 7972 1517 7987 1523
rect 4237 1497 4275 1503
rect 4356 1497 4387 1503
rect 4404 1497 4419 1503
rect 5517 1497 5539 1503
rect 5597 1497 5651 1503
rect 6116 1497 6131 1503
rect 6308 1497 6323 1503
rect 6333 1497 6435 1503
rect 6660 1497 6675 1503
rect 6916 1497 6931 1503
rect 7069 1497 7084 1503
rect 7165 1497 7180 1503
rect 7204 1497 7219 1503
rect 7597 1497 7619 1503
rect 301 1477 332 1483
rect 381 1477 412 1483
rect 548 1477 563 1483
rect 1412 1477 1427 1483
rect 1453 1477 1507 1483
rect 1700 1477 1731 1483
rect 1757 1477 1859 1483
rect 2564 1477 2579 1483
rect 3277 1477 3347 1483
rect 3581 1477 3628 1483
rect 4068 1477 4083 1483
rect 4324 1477 4339 1483
rect 4349 1477 4364 1483
rect 5197 1477 5219 1483
rect 6045 1477 6067 1483
rect 6349 1477 6380 1483
rect 6477 1477 6499 1483
rect 6765 1477 6780 1483
rect 6893 1477 6947 1483
rect 6973 1477 6988 1483
rect 7021 1477 7043 1483
rect 8109 1477 8156 1483
rect 4620 1464 4628 1472
rect 3709 1457 3756 1463
rect 5308 1463 5316 1472
rect 5308 1457 5340 1463
rect 356 1436 358 1444
rect 500 1436 502 1444
rect 1549 1437 1564 1443
rect 2196 1436 2198 1444
rect 8052 1436 8056 1444
rect 3272 1406 3278 1414
rect 3286 1406 3292 1414
rect 3300 1406 3306 1414
rect 3314 1406 3320 1414
rect 6344 1406 6350 1414
rect 6358 1406 6364 1414
rect 6372 1406 6378 1414
rect 6386 1406 6392 1414
rect 522 1376 524 1384
rect 1258 1376 1260 1384
rect 1306 1376 1308 1384
rect 2138 1376 2140 1384
rect 5384 1376 5388 1384
rect 5677 1377 5692 1383
rect 6120 1376 6124 1384
rect 7764 1377 7779 1383
rect 541 1337 556 1343
rect 2221 1337 2275 1343
rect 2381 1337 2435 1343
rect 2717 1337 2739 1343
rect 3789 1337 3811 1343
rect 3997 1343 4003 1363
rect 4445 1357 4467 1363
rect 5284 1357 5299 1363
rect 3997 1337 4012 1343
rect 4404 1337 4419 1343
rect 4557 1337 4579 1343
rect 5261 1337 5276 1343
rect 5421 1337 5436 1343
rect 6045 1337 6067 1343
rect 6605 1337 6659 1343
rect 7636 1337 7651 1343
rect 7933 1337 7948 1343
rect 477 1317 515 1323
rect 621 1317 643 1323
rect 653 1317 668 1323
rect 509 1297 515 1317
rect 1213 1317 1251 1323
rect 1357 1317 1372 1323
rect 1245 1297 1251 1317
rect 1405 1317 1436 1323
rect 2013 1317 2051 1323
rect 2084 1317 2099 1323
rect 2285 1317 2332 1323
rect 2477 1317 2500 1323
rect 2492 1314 2500 1317
rect 3364 1317 3427 1323
rect 3437 1317 3491 1323
rect 3613 1317 3628 1323
rect 3773 1317 3788 1323
rect 3949 1317 3964 1323
rect 4388 1317 4403 1323
rect 4493 1317 4547 1323
rect 4685 1317 4716 1323
rect 4797 1317 4860 1323
rect 5204 1317 5219 1323
rect 5821 1317 5843 1323
rect 5901 1317 5923 1323
rect 6004 1317 6019 1323
rect 6493 1317 6531 1323
rect 1357 1297 1379 1303
rect 1396 1296 1404 1304
rect 2068 1297 2083 1303
rect 4356 1296 4364 1304
rect 6525 1297 6531 1317
rect 7565 1317 7619 1323
rect 7677 1317 7731 1323
rect 1292 1283 1300 1288
rect 1532 1284 1540 1288
rect 2124 1284 2132 1288
rect 1284 1277 1300 1283
rect 1466 1276 1468 1284
rect 4173 1277 4220 1283
rect 4173 1257 4179 1277
rect 4564 1277 4579 1283
rect 7725 1277 7772 1283
rect 4292 1256 4294 1264
rect 3341 1237 3388 1243
rect 4746 1236 4748 1244
rect 4938 1236 4940 1244
rect 6554 1236 6556 1244
rect 6932 1236 6934 1244
rect 1736 1206 1742 1214
rect 1750 1206 1756 1214
rect 1764 1206 1770 1214
rect 1778 1206 1784 1214
rect 4808 1206 4814 1214
rect 4822 1206 4828 1214
rect 4836 1206 4842 1214
rect 4850 1206 4856 1214
rect 3434 1176 3436 1184
rect 5220 1176 5222 1184
rect 7242 1176 7244 1184
rect 7338 1176 7340 1184
rect 5338 1156 5340 1164
rect 868 1136 870 1144
rect 2618 1136 2620 1144
rect 6756 1137 6787 1143
rect 8140 1137 8156 1143
rect 6620 1132 6628 1136
rect 8140 1132 8148 1137
rect 541 1097 556 1103
rect 580 1097 595 1103
rect 829 1103 835 1123
rect 829 1097 860 1103
rect 893 1103 899 1123
rect 996 1117 1011 1123
rect 893 1097 931 1103
rect 1053 1097 1075 1103
rect 1229 1103 1235 1123
rect 1181 1097 1219 1103
rect 1229 1097 1267 1103
rect 1725 1103 1731 1123
rect 1693 1097 1731 1103
rect 2029 1097 2051 1103
rect 2212 1097 2243 1103
rect 2420 1097 2435 1103
rect 2508 1103 2516 1108
rect 2508 1097 2531 1103
rect 1044 1077 1059 1083
rect 1085 1077 1139 1083
rect 1501 1077 1523 1083
rect 1501 1064 1507 1077
rect 1764 1077 1804 1083
rect 2125 1077 2140 1083
rect 2525 1077 2531 1097
rect 2589 1103 2595 1123
rect 4740 1116 4748 1124
rect 4916 1117 4931 1123
rect 4948 1116 4956 1124
rect 5149 1117 5171 1123
rect 5300 1117 5315 1123
rect 5837 1117 5868 1123
rect 6260 1116 6268 1124
rect 2557 1097 2595 1103
rect 2749 1097 2771 1103
rect 3613 1097 3651 1103
rect 3668 1097 3683 1103
rect 4148 1097 4163 1103
rect 4173 1097 4227 1103
rect 4989 1103 4995 1116
rect 4772 1097 4787 1103
rect 4957 1097 4995 1103
rect 5252 1097 5283 1103
rect 5540 1097 5555 1103
rect 5716 1097 5747 1103
rect 5805 1097 5843 1103
rect 6141 1097 6156 1103
rect 6660 1097 6691 1103
rect 7341 1097 7379 1103
rect 2845 1077 2867 1083
rect 3236 1077 3251 1083
rect 3460 1077 3491 1083
rect 3517 1077 3571 1083
rect 4100 1077 4115 1083
rect 4125 1077 4140 1083
rect 2477 1057 2492 1063
rect 4109 1057 4115 1077
rect 7373 1084 7379 1097
rect 7629 1103 7635 1123
rect 7693 1117 7731 1123
rect 8093 1117 8131 1123
rect 7533 1097 7587 1103
rect 7597 1097 7635 1103
rect 7668 1097 7699 1103
rect 7805 1097 7843 1103
rect 7917 1097 7932 1103
rect 8045 1097 8083 1103
rect 4973 1077 4988 1083
rect 5165 1077 5203 1083
rect 5416 1076 5420 1084
rect 5645 1077 5667 1083
rect 5853 1077 5875 1083
rect 5885 1077 5916 1083
rect 5853 1064 5859 1077
rect 5956 1077 5971 1083
rect 6077 1077 6131 1083
rect 6285 1077 6307 1083
rect 6628 1077 6643 1083
rect 6653 1077 6668 1083
rect 7156 1077 7171 1083
rect 7261 1077 7299 1083
rect 7405 1077 7420 1083
rect 7949 1077 8003 1083
rect 6669 1057 6675 1076
rect 244 1036 248 1044
rect 820 1036 822 1044
rect 1140 1036 1142 1044
rect 1428 1036 1430 1044
rect 1540 1036 1542 1044
rect 1604 1036 1608 1044
rect 1738 1036 1740 1044
rect 4820 1037 4867 1043
rect 8004 1036 8006 1044
rect 3272 1006 3278 1014
rect 3286 1006 3292 1014
rect 3300 1006 3306 1014
rect 3314 1006 3320 1014
rect 6344 1006 6350 1014
rect 6358 1006 6364 1014
rect 6372 1006 6378 1014
rect 6386 1006 6392 1014
rect 788 977 803 983
rect 3636 976 3638 984
rect 4376 976 4380 984
rect 4874 976 4876 984
rect 5636 976 5638 984
rect 7034 976 7036 984
rect 429 957 451 963
rect 4125 957 4147 963
rect 6637 957 6659 963
rect 7101 957 7124 963
rect 7116 954 7124 957
rect 7644 944 7652 954
rect 845 937 899 943
rect 925 937 956 943
rect 1629 937 1683 943
rect 2724 937 2740 943
rect 3076 937 3091 943
rect 3236 937 3251 943
rect 3501 937 3523 943
rect 4493 937 4547 943
rect 4573 937 4588 943
rect 4797 937 4860 943
rect 4957 937 5011 943
rect 5709 937 5731 943
rect 6189 937 6204 943
rect 6221 937 6259 943
rect 6333 937 6380 943
rect 7037 937 7091 943
rect 7384 937 7404 943
rect 7821 937 7843 943
rect 212 917 227 923
rect 285 917 300 923
rect 349 917 364 923
rect 452 917 467 923
rect 477 917 499 923
rect 605 917 627 923
rect 989 917 1027 923
rect 221 897 259 903
rect 1021 897 1027 917
rect 1053 917 1107 923
rect 1124 917 1155 923
rect 2493 917 2515 923
rect 2557 917 2595 923
rect 1197 897 1228 903
rect 1252 896 1260 904
rect 2589 897 2595 917
rect 2644 917 2659 923
rect 2669 917 2684 923
rect 2941 917 2972 923
rect 2989 917 3027 923
rect 3021 897 3027 917
rect 3101 917 3155 923
rect 3277 917 3292 923
rect 3741 917 3779 923
rect 3741 897 3747 917
rect 3981 917 4019 923
rect 4013 897 4019 917
rect 4148 917 4163 923
rect 4173 917 4195 923
rect 4253 917 4268 923
rect 4589 917 4627 923
rect 4637 917 4675 923
rect 4637 897 4643 917
rect 5181 917 5203 923
rect 5693 917 5708 923
rect 6413 917 6435 923
rect 6637 917 6652 923
rect 6957 917 6995 923
rect 7437 923 7443 936
rect 7420 917 7443 923
rect 7420 912 7428 917
rect 6164 896 6172 904
rect 7412 897 7427 903
rect 7533 897 7548 903
rect 7860 896 7868 904
rect 282 876 284 884
rect 346 876 348 884
rect 621 877 636 883
rect 692 876 696 884
rect 1764 877 1795 883
rect 3300 877 3372 883
rect 3444 876 3448 884
rect 4042 876 4044 884
rect 4860 883 4868 888
rect 4852 877 4868 883
rect 5028 877 5043 883
rect 6536 876 6540 884
rect 1508 836 1510 844
rect 2484 836 2486 844
rect 3050 836 3052 844
rect 4778 836 4780 844
rect 7338 836 7340 844
rect 1736 806 1742 814
rect 1750 806 1756 814
rect 1764 806 1770 814
rect 1778 806 1784 814
rect 4808 806 4814 814
rect 4822 806 4828 814
rect 4836 806 4842 814
rect 4850 806 4856 814
rect 1338 776 1340 784
rect 4116 776 4118 784
rect 1236 737 1252 743
rect 1244 732 1252 737
rect 1380 737 1411 743
rect 5562 736 5564 744
rect 7180 732 7188 736
rect 77 703 83 723
rect 45 697 83 703
rect 109 697 163 703
rect 180 697 195 703
rect 893 697 908 703
rect 1085 697 1116 703
rect 1309 697 1331 703
rect 2301 703 2307 723
rect 2324 716 2332 724
rect 2525 717 2547 723
rect 5108 716 5116 724
rect 3612 706 3620 716
rect 2269 697 2307 703
rect 2484 697 2515 703
rect 2612 697 2627 703
rect 2813 697 2844 703
rect 2884 697 2899 703
rect 3044 697 3059 703
rect 3396 697 3411 703
rect 3421 697 3443 703
rect 3892 697 3923 703
rect 4020 696 4024 704
rect 4148 697 4179 703
rect 5133 703 5139 723
rect 5133 697 5155 703
rect 5469 697 5491 703
rect 5420 692 5428 696
rect 205 677 220 683
rect 205 657 211 677
rect 237 677 252 683
rect 404 677 420 683
rect 1124 676 1126 684
rect 1277 677 1292 683
rect 1517 677 1539 683
rect 1613 677 1667 683
rect 1821 677 1843 683
rect 2541 677 2556 683
rect 2628 677 2643 683
rect 2861 677 2883 683
rect 4196 677 4211 683
rect 5156 677 5171 683
rect 5485 684 5491 697
rect 5700 697 5715 703
rect 5965 703 5971 723
rect 5917 697 5955 703
rect 5965 697 6003 703
rect 6525 703 6531 723
rect 7604 716 7608 724
rect 8116 716 8124 724
rect 8141 717 8156 723
rect 6020 697 6035 703
rect 6525 697 6563 703
rect 6733 697 6771 703
rect 7197 697 7235 703
rect 7469 697 7507 703
rect 7693 697 7715 703
rect 6340 677 6403 683
rect 6573 677 6595 683
rect 1357 657 1379 663
rect 2012 663 2020 672
rect 6589 664 6595 677
rect 7293 677 7315 683
rect 7380 677 7395 683
rect 7556 677 7571 683
rect 7661 677 7676 683
rect 7821 677 7836 683
rect 1988 657 2020 663
rect 3373 657 3395 663
rect 6045 657 6060 663
rect 356 636 358 644
rect 1396 637 1411 643
rect 6468 636 6470 644
rect 6516 636 6518 644
rect 7928 636 7932 644
rect 3272 606 3278 614
rect 3286 606 3292 614
rect 3300 606 3306 614
rect 3314 606 3320 614
rect 6344 606 6350 614
rect 6358 606 6364 614
rect 6372 606 6378 614
rect 6386 606 6392 614
rect 2184 576 2188 584
rect 2376 576 2380 584
rect 2676 576 2678 584
rect 2868 576 2870 584
rect 317 557 332 563
rect 1556 556 1564 564
rect 4829 557 4892 563
rect 4973 557 4988 563
rect 7884 557 7907 563
rect 7981 557 8003 563
rect 221 537 252 543
rect 349 537 403 543
rect 541 537 563 543
rect 909 537 924 543
rect 1949 537 1971 543
rect 2237 543 2243 556
rect 7884 554 7892 557
rect 2221 537 2243 543
rect 3661 537 3683 543
rect 4141 537 4163 543
rect 4588 537 4612 543
rect 5069 537 5123 543
rect 5485 537 5507 543
rect 5645 537 5699 543
rect 6173 537 6220 543
rect 6445 537 6460 543
rect 7692 537 7716 543
rect 7940 537 7955 543
rect 8045 537 8060 543
rect 100 517 131 523
rect 237 517 275 523
rect 301 517 339 523
rect 237 497 243 517
rect 1133 517 1148 523
rect 1277 517 1299 523
rect 1565 517 1603 523
rect 1613 517 1644 523
rect 1565 504 1571 517
rect 2797 517 2835 523
rect 3149 517 3171 523
rect 3325 517 3340 523
rect 4317 517 4371 523
rect 4516 517 4531 523
rect 5181 523 5187 536
rect 5165 517 5187 523
rect 5197 517 5235 523
rect 516 496 524 504
rect 4253 497 4268 503
rect 5229 497 5235 517
rect 5549 517 5587 523
rect 5549 497 5555 517
rect 5757 517 5788 523
rect 5972 517 5987 523
rect 6109 517 6147 523
rect 6109 497 6115 517
rect 6541 517 6595 523
rect 6605 517 6643 523
rect 6637 497 6643 517
rect 6781 517 6835 523
rect 6868 517 6899 523
rect 6909 517 6931 523
rect 7101 517 7155 523
rect 7181 517 7219 523
rect 7229 517 7251 523
rect 6861 497 6867 516
rect 7181 504 7187 517
rect 7364 517 7395 523
rect 7917 517 7939 523
rect 7468 484 7476 488
rect 1628 477 1644 483
rect 1700 477 1747 483
rect 2797 477 2812 483
rect 6666 476 6668 484
rect 6973 477 6988 483
rect 8068 477 8083 483
rect 1306 436 1308 444
rect 3178 436 3180 444
rect 7156 436 7158 444
rect 1736 406 1742 414
rect 1750 406 1756 414
rect 1764 406 1770 414
rect 1778 406 1784 414
rect 4808 406 4814 414
rect 4822 406 4828 414
rect 4836 406 4842 414
rect 4850 406 4856 414
rect 628 337 643 343
rect 1738 336 1740 344
rect 3556 336 3558 344
rect 5066 336 5068 344
rect 5597 343 5603 363
rect 5597 337 5644 343
rect 5748 336 5750 344
rect 1629 317 1651 323
rect 1668 316 1676 324
rect 404 297 419 303
rect 1181 297 1219 303
rect 1229 297 1244 303
rect 1885 284 1891 303
rect 2445 297 2467 303
rect 2717 303 2723 323
rect 2740 316 2748 324
rect 2820 317 2835 323
rect 3300 317 3331 323
rect 3469 317 3484 323
rect 2685 297 2723 303
rect 3517 303 3523 323
rect 3492 297 3507 303
rect 3517 297 3548 303
rect 3581 303 3587 323
rect 3940 316 3948 324
rect 3581 297 3619 303
rect 3965 303 3971 323
rect 3924 297 3939 303
rect 3965 297 3987 303
rect 4413 297 4428 303
rect 4484 297 4499 303
rect 4909 297 4931 303
rect 5037 303 5043 323
rect 5204 317 5219 323
rect 5812 316 5820 324
rect 6845 317 6883 323
rect 5005 297 5043 303
rect 5405 297 5427 303
rect 909 277 931 283
rect 1812 277 1843 283
rect 1892 277 1907 283
rect 2349 277 2371 283
rect 2644 277 2659 283
rect 2872 276 2876 284
rect 2973 277 3027 283
rect 3437 277 3475 283
rect 3741 277 3756 283
rect 1100 263 1108 272
rect 1076 257 1108 263
rect 2316 263 2324 266
rect 3741 264 3747 277
rect 3837 277 3859 283
rect 3988 277 4003 283
rect 4349 277 4403 283
rect 4477 277 4492 283
rect 5405 277 5411 297
rect 5501 297 5523 303
rect 5533 297 5548 303
rect 5693 297 5747 303
rect 5796 297 5811 303
rect 5885 297 5939 303
rect 7748 297 7779 303
rect 8100 297 8115 303
rect 6093 277 6108 283
rect 6301 277 6323 283
rect 6900 277 6915 283
rect 7613 277 7651 283
rect 7716 277 7731 283
rect 7917 283 7923 296
rect 7901 277 7923 283
rect 8141 277 8156 283
rect 2316 257 2339 263
rect 4932 257 4947 263
rect 602 236 604 244
rect 1304 236 1308 244
rect 2794 236 2796 244
rect 4792 236 4796 244
rect 5178 236 5180 244
rect 5348 236 5352 244
rect 6836 236 6838 244
rect 3272 206 3278 214
rect 3286 206 3292 214
rect 3300 206 3306 214
rect 3314 206 3320 214
rect 6344 206 6350 214
rect 6358 206 6364 214
rect 6372 206 6378 214
rect 6386 206 6392 214
rect 292 176 294 184
rect 552 176 556 184
rect 714 176 716 184
rect 1162 176 1164 184
rect 1757 177 1804 183
rect 2548 176 2550 184
rect 2826 176 2828 184
rect 4026 176 4028 184
rect 4372 176 4374 184
rect 4490 176 4492 184
rect 8100 177 8115 183
rect 173 143 179 163
rect 1437 157 1459 163
rect 1652 156 1660 164
rect 3764 156 3772 164
rect 4813 157 4844 163
rect 7101 157 7124 163
rect 164 137 179 143
rect 260 137 275 143
rect 333 137 387 143
rect 596 137 611 143
rect 676 137 691 143
rect 1132 137 1148 143
rect 1396 137 1411 143
rect 3949 143 3955 156
rect 7116 154 7124 157
rect 7500 157 7532 163
rect 7500 148 7508 157
rect 3949 137 3971 143
rect 4868 137 4899 143
rect 5268 137 5283 143
rect 6541 137 6563 143
rect 6852 137 6867 143
rect 6884 137 6899 143
rect 6909 137 6963 143
rect 7069 137 7091 143
rect 7325 137 7363 143
rect 7644 137 7668 143
rect 356 117 371 123
rect 861 117 915 123
rect 1021 117 1036 123
rect 1060 117 1075 123
rect 1485 117 1516 123
rect 1876 117 1891 123
rect 2093 117 2147 123
rect 2196 117 2211 123
rect 2877 117 2908 123
rect 2941 117 2979 123
rect 93 97 115 103
rect 1597 97 1612 103
rect 1629 97 1651 103
rect 2260 97 2275 103
rect 2676 96 2680 104
rect 2852 97 2867 103
rect 2973 97 2979 117
rect 3140 117 3155 123
rect 3981 117 4019 123
rect 3677 97 3692 103
rect 4013 97 4019 117
rect 5964 124 5972 128
rect 4381 117 4419 123
rect 4381 97 4387 117
rect 4621 117 4659 123
rect 4653 97 4659 117
rect 4692 117 4723 123
rect 4733 117 4787 123
rect 4717 97 4723 117
rect 5245 117 5267 123
rect 5476 117 5491 123
rect 6509 117 6524 123
rect 6701 117 6755 123
rect 6877 117 6892 123
rect 7901 117 7932 123
rect 7044 96 7052 104
rect 7341 97 7356 103
rect 7428 96 7436 104
rect 138 76 140 84
rect 772 76 774 84
rect 1892 76 1894 84
rect 1949 77 1964 83
rect 5656 76 5660 84
rect 7452 77 7475 83
rect 1736 6 1742 14
rect 1750 6 1756 14
rect 1764 6 1770 14
rect 1778 6 1784 14
rect 4808 6 4814 14
rect 4822 6 4828 14
rect 4836 6 4842 14
rect 4850 6 4856 14
<< m2contact >>
rect 3278 5806 3286 5814
rect 3292 5806 3300 5814
rect 3306 5806 3314 5814
rect 6350 5806 6358 5814
rect 6364 5806 6372 5814
rect 6378 5806 6386 5814
rect 2364 5776 2372 5784
rect 2828 5776 2836 5784
rect 3292 5776 3300 5784
rect 3660 5776 3668 5784
rect 3932 5776 3940 5784
rect 4172 5776 4180 5784
rect 4764 5776 4772 5784
rect 5036 5776 5044 5784
rect 6204 5776 6212 5784
rect 284 5756 292 5764
rect 428 5756 436 5764
rect 636 5756 644 5764
rect 940 5756 948 5764
rect 1036 5756 1044 5764
rect 1068 5756 1076 5764
rect 1276 5756 1284 5764
rect 1484 5756 1492 5764
rect 1868 5756 1876 5764
rect 2460 5756 2468 5764
rect 2732 5756 2740 5764
rect 3148 5756 3156 5764
rect 3676 5756 3684 5764
rect 4156 5756 4164 5764
rect 4380 5756 4388 5764
rect 4556 5756 4564 5764
rect 4780 5756 4788 5764
rect 5052 5756 5060 5764
rect 5580 5756 5588 5764
rect 5612 5756 5620 5764
rect 5676 5756 5684 5764
rect 5740 5756 5748 5764
rect 5836 5756 5844 5764
rect 6140 5756 6148 5764
rect 6188 5756 6196 5764
rect 7164 5756 7172 5764
rect 332 5732 340 5740
rect 364 5736 372 5744
rect 860 5736 868 5744
rect 876 5736 884 5744
rect 972 5736 980 5744
rect 1148 5736 1156 5744
rect 1260 5736 1268 5744
rect 1324 5736 1332 5744
rect 1692 5736 1700 5744
rect 1836 5736 1844 5744
rect 1980 5736 1988 5744
rect 2012 5736 2020 5744
rect 2204 5736 2212 5744
rect 2508 5736 2516 5744
rect 2540 5736 2548 5744
rect 2572 5736 2580 5744
rect 2604 5736 2612 5744
rect 2668 5736 2676 5744
rect 2700 5736 2708 5744
rect 2988 5736 2996 5744
rect 3020 5736 3028 5744
rect 3084 5736 3092 5744
rect 3116 5736 3124 5744
rect 3452 5736 3460 5744
rect 3740 5736 3748 5744
rect 3804 5736 3812 5744
rect 3836 5736 3844 5744
rect 3868 5736 3876 5744
rect 3964 5736 3972 5744
rect 3996 5736 4004 5744
rect 4028 5736 4036 5744
rect 4332 5736 4340 5744
rect 4396 5736 4404 5744
rect 4492 5736 4500 5744
rect 4524 5736 4532 5744
rect 4972 5736 4980 5744
rect 4988 5736 4996 5744
rect 5084 5736 5092 5744
rect 5132 5736 5140 5744
rect 5180 5736 5188 5744
rect 5212 5736 5220 5744
rect 5388 5736 5396 5744
rect 5452 5736 5460 5744
rect 5484 5736 5492 5744
rect 5500 5736 5508 5744
rect 5564 5736 5572 5744
rect 5612 5736 5620 5744
rect 5708 5736 5716 5744
rect 5852 5736 5860 5744
rect 5884 5736 5892 5744
rect 5900 5736 5908 5744
rect 5916 5736 5924 5744
rect 5948 5736 5956 5744
rect 6044 5736 6052 5744
rect 6364 5736 6372 5744
rect 6444 5736 6452 5744
rect 6572 5736 6580 5744
rect 6780 5736 6788 5744
rect 7052 5736 7060 5744
rect 7116 5736 7124 5744
rect 7148 5736 7156 5744
rect 7196 5736 7204 5744
rect 7228 5736 7236 5744
rect 7324 5736 7332 5744
rect 7340 5736 7348 5744
rect 7436 5736 7444 5744
rect 7612 5736 7620 5744
rect 7692 5736 7700 5744
rect 7836 5736 7844 5744
rect 7964 5736 7972 5744
rect 7996 5736 8004 5744
rect 92 5716 100 5724
rect 124 5716 132 5724
rect 204 5716 212 5724
rect 236 5716 244 5724
rect 380 5716 388 5724
rect 508 5716 516 5724
rect 556 5716 564 5724
rect 684 5716 692 5724
rect 700 5716 708 5724
rect 924 5716 932 5724
rect 988 5716 996 5724
rect 1004 5716 1012 5724
rect 1036 5716 1044 5724
rect 1116 5716 1124 5724
rect 1164 5716 1172 5724
rect 204 5696 212 5704
rect 396 5696 404 5704
rect 716 5696 724 5704
rect 908 5696 916 5704
rect 1132 5696 1140 5704
rect 1196 5696 1204 5704
rect 1244 5716 1252 5724
rect 1340 5716 1348 5724
rect 1420 5718 1428 5726
rect 1484 5716 1492 5724
rect 1596 5716 1604 5724
rect 1644 5716 1652 5724
rect 1676 5716 1684 5724
rect 1788 5716 1796 5724
rect 1820 5716 1828 5724
rect 2060 5716 2068 5724
rect 2268 5716 2276 5724
rect 2284 5716 2292 5724
rect 2380 5716 2388 5724
rect 2412 5716 2420 5724
rect 2588 5716 2596 5724
rect 2652 5716 2660 5724
rect 2732 5716 2740 5724
rect 2780 5716 2788 5724
rect 2812 5716 2820 5724
rect 2924 5716 2932 5724
rect 3068 5716 3076 5724
rect 3148 5716 3156 5724
rect 3196 5716 3204 5724
rect 3276 5716 3284 5724
rect 3356 5716 3364 5724
rect 3404 5716 3412 5724
rect 3548 5716 3556 5724
rect 3596 5716 3604 5724
rect 3724 5716 3732 5724
rect 1276 5696 1284 5704
rect 1356 5696 1364 5704
rect 1612 5696 1620 5704
rect 1628 5696 1636 5704
rect 1724 5696 1732 5704
rect 1788 5696 1796 5704
rect 2380 5696 2388 5704
rect 2476 5696 2484 5704
rect 2492 5696 2500 5704
rect 2620 5696 2628 5704
rect 2636 5696 2644 5704
rect 2812 5696 2820 5704
rect 3036 5696 3044 5704
rect 3052 5696 3060 5704
rect 3228 5696 3236 5704
rect 3884 5716 3892 5724
rect 3900 5716 3908 5724
rect 3948 5716 3956 5724
rect 3772 5696 3780 5704
rect 4060 5696 4068 5704
rect 4092 5716 4100 5724
rect 4108 5716 4116 5724
rect 4284 5716 4292 5724
rect 4460 5716 4468 5724
rect 4508 5716 4516 5724
rect 4556 5716 4564 5724
rect 4620 5718 4628 5726
rect 4684 5716 4692 5724
rect 4844 5716 4852 5724
rect 5004 5716 5012 5724
rect 5068 5716 5076 5724
rect 5244 5718 5252 5726
rect 5612 5716 5620 5724
rect 5692 5716 5700 5724
rect 5788 5716 5796 5724
rect 5868 5716 5876 5724
rect 5932 5716 5940 5724
rect 5980 5716 5988 5724
rect 6076 5716 6084 5724
rect 6092 5716 6100 5724
rect 6156 5716 6164 5724
rect 6316 5716 6324 5724
rect 6652 5716 6660 5724
rect 6716 5718 6724 5726
rect 6956 5716 6964 5724
rect 7004 5716 7012 5724
rect 7020 5716 7028 5724
rect 7100 5716 7108 5724
rect 7132 5716 7140 5724
rect 7212 5716 7220 5724
rect 7580 5718 7588 5726
rect 7708 5716 7716 5724
rect 8028 5718 8036 5726
rect 5116 5696 5124 5704
rect 5180 5696 5188 5704
rect 5420 5696 5428 5704
rect 5516 5696 5524 5704
rect 5660 5696 5668 5704
rect 5804 5696 5812 5704
rect 5820 5696 5828 5704
rect 6060 5696 6068 5704
rect 6972 5696 6980 5704
rect 6988 5696 6996 5704
rect 7084 5696 7092 5704
rect 7100 5696 7108 5704
rect 7260 5696 7268 5704
rect 636 5676 644 5684
rect 1100 5676 1108 5684
rect 1244 5676 1252 5684
rect 1324 5676 1332 5684
rect 1516 5676 1524 5684
rect 1580 5676 1588 5684
rect 4204 5676 4212 5684
rect 5340 5676 5348 5684
rect 5372 5676 5380 5684
rect 5484 5676 5492 5684
rect 5772 5676 5780 5684
rect 6940 5676 6948 5684
rect 1116 5656 1124 5664
rect 188 5636 196 5644
rect 300 5636 308 5644
rect 412 5636 420 5644
rect 748 5636 756 5644
rect 1004 5636 1012 5644
rect 1548 5636 1556 5644
rect 1564 5636 1572 5644
rect 1820 5636 1828 5644
rect 2172 5636 2180 5644
rect 2540 5636 2548 5644
rect 2668 5636 2676 5644
rect 3084 5636 3092 5644
rect 3836 5636 3844 5644
rect 3996 5636 4004 5644
rect 4364 5636 4372 5644
rect 4748 5636 4756 5644
rect 5740 5636 5748 5644
rect 5788 5636 5796 5644
rect 6204 5636 6212 5644
rect 6588 5636 6596 5644
rect 6892 5636 6900 5644
rect 6956 5636 6964 5644
rect 7164 5636 7172 5644
rect 7404 5636 7412 5644
rect 7452 5636 7460 5644
rect 7820 5636 7828 5644
rect 8156 5636 8164 5644
rect 1742 5606 1750 5614
rect 1756 5606 1764 5614
rect 1770 5606 1778 5614
rect 4814 5606 4822 5614
rect 4828 5606 4836 5614
rect 4842 5606 4850 5614
rect 364 5576 372 5584
rect 492 5576 500 5584
rect 956 5576 964 5584
rect 1020 5576 1028 5584
rect 1884 5576 1892 5584
rect 1980 5576 1988 5584
rect 2252 5576 2260 5584
rect 2332 5576 2340 5584
rect 2444 5576 2452 5584
rect 4108 5576 4116 5584
rect 4172 5576 4180 5584
rect 4492 5576 4500 5584
rect 4620 5576 4628 5584
rect 5468 5576 5476 5584
rect 5532 5576 5540 5584
rect 5740 5576 5748 5584
rect 5996 5576 6004 5584
rect 6092 5576 6100 5584
rect 6748 5576 6756 5584
rect 7132 5576 7140 5584
rect 7212 5576 7220 5584
rect 7276 5576 7284 5584
rect 7324 5576 7332 5584
rect 556 5556 564 5564
rect 1244 5556 1252 5564
rect 1932 5556 1940 5564
rect 4380 5556 4388 5564
rect 4556 5556 4564 5564
rect 4812 5556 4820 5564
rect 5900 5556 5908 5564
rect 7868 5556 7876 5564
rect 7948 5556 7956 5564
rect 492 5536 500 5544
rect 572 5536 580 5544
rect 1468 5536 1476 5544
rect 1996 5536 2004 5544
rect 2028 5536 2036 5544
rect 2172 5536 2180 5544
rect 4572 5536 4580 5544
rect 5020 5536 5028 5544
rect 5100 5536 5108 5544
rect 5164 5536 5172 5544
rect 5772 5536 5780 5544
rect 5836 5536 5844 5544
rect 7084 5536 7092 5544
rect 7148 5536 7156 5544
rect 7340 5536 7348 5544
rect 7884 5536 7892 5544
rect 7996 5536 8004 5544
rect 332 5516 340 5524
rect 396 5516 404 5524
rect 476 5516 484 5524
rect 540 5516 548 5524
rect 76 5496 84 5504
rect 124 5496 132 5504
rect 204 5496 212 5504
rect 268 5496 276 5504
rect 284 5496 292 5504
rect 364 5496 372 5504
rect 428 5496 436 5504
rect 508 5496 516 5504
rect 556 5496 564 5504
rect 748 5496 756 5504
rect 796 5496 804 5504
rect 972 5496 980 5504
rect 1036 5496 1044 5504
rect 1052 5496 1060 5504
rect 1100 5516 1108 5524
rect 1148 5516 1156 5524
rect 1340 5516 1348 5524
rect 1404 5516 1412 5524
rect 1180 5496 1188 5504
rect 1356 5496 1364 5504
rect 1372 5496 1380 5504
rect 1436 5496 1444 5504
rect 1964 5516 1972 5524
rect 2204 5516 2212 5524
rect 2220 5516 2228 5524
rect 2636 5516 2644 5524
rect 2860 5516 2868 5524
rect 2908 5516 2916 5524
rect 3148 5516 3156 5524
rect 3436 5516 3444 5524
rect 3532 5516 3540 5524
rect 3548 5516 3556 5524
rect 4044 5516 4052 5524
rect 4220 5516 4228 5524
rect 4332 5516 4340 5524
rect 4348 5516 4356 5524
rect 4412 5516 4420 5524
rect 4524 5516 4532 5524
rect 4540 5516 4548 5524
rect 4780 5516 4788 5524
rect 4924 5516 4932 5524
rect 4940 5516 4948 5524
rect 4972 5516 4980 5524
rect 5004 5516 5012 5524
rect 5068 5516 5076 5524
rect 5132 5516 5140 5524
rect 5516 5516 5524 5524
rect 5804 5516 5812 5524
rect 5868 5516 5876 5524
rect 6028 5516 6036 5524
rect 6140 5516 6148 5524
rect 6684 5516 6692 5524
rect 6780 5516 6788 5524
rect 7116 5516 7124 5524
rect 7596 5516 7604 5524
rect 7852 5516 7860 5524
rect 7916 5516 7924 5524
rect 8076 5516 8084 5524
rect 1612 5494 1620 5502
rect 1660 5496 1668 5504
rect 1852 5496 1860 5504
rect 1932 5496 1940 5504
rect 1980 5496 1988 5504
rect 2092 5496 2100 5504
rect 2156 5496 2164 5504
rect 2220 5496 2228 5504
rect 2252 5496 2260 5504
rect 2428 5496 2436 5504
rect 2476 5496 2484 5504
rect 2716 5496 2724 5504
rect 2764 5496 2772 5504
rect 2844 5496 2852 5504
rect 2940 5496 2948 5504
rect 3004 5494 3012 5502
rect 3324 5496 3332 5504
rect 3356 5496 3364 5504
rect 3436 5496 3444 5504
rect 3468 5496 3476 5504
rect 3580 5496 3588 5504
rect 3644 5496 3652 5504
rect 3708 5494 3716 5502
rect 3772 5496 3780 5504
rect 3916 5496 3924 5504
rect 3980 5494 3988 5502
rect 4044 5496 4052 5504
rect 4124 5496 4132 5504
rect 4380 5496 4388 5504
rect 4444 5496 4452 5504
rect 220 5476 228 5484
rect 252 5476 260 5484
rect 300 5476 308 5484
rect 380 5476 388 5484
rect 604 5476 612 5484
rect 844 5476 852 5484
rect 876 5476 884 5484
rect 892 5480 900 5488
rect 988 5476 996 5484
rect 1020 5476 1028 5484
rect 1052 5476 1060 5484
rect 1132 5476 1140 5484
rect 1196 5476 1204 5484
rect 1276 5480 1284 5488
rect 1292 5476 1300 5484
rect 1308 5476 1316 5484
rect 1340 5476 1348 5484
rect 1388 5476 1396 5484
rect 1420 5476 1428 5484
rect 1452 5476 1460 5484
rect 1836 5476 1844 5484
rect 1948 5476 1956 5484
rect 2092 5476 2100 5484
rect 2108 5476 2116 5484
rect 2172 5476 2180 5484
rect 2444 5476 2452 5484
rect 2492 5476 2500 5484
rect 2668 5476 2676 5484
rect 2700 5476 2708 5484
rect 2796 5476 2804 5484
rect 2828 5476 2836 5484
rect 2892 5476 2900 5484
rect 2940 5476 2948 5484
rect 3212 5476 3220 5484
rect 3564 5476 3572 5484
rect 3596 5476 3604 5484
rect 3628 5476 3636 5484
rect 3676 5476 3684 5484
rect 4012 5476 4020 5484
rect 4076 5476 4084 5484
rect 4252 5476 4260 5484
rect 4268 5476 4276 5484
rect 4396 5476 4404 5484
rect 4460 5476 4468 5484
rect 4492 5496 4500 5504
rect 4556 5496 4564 5504
rect 4780 5496 4788 5504
rect 4972 5496 4980 5504
rect 5020 5496 5028 5504
rect 5068 5496 5076 5504
rect 5100 5496 5108 5504
rect 5148 5496 5156 5504
rect 5180 5496 5188 5504
rect 5260 5496 5268 5504
rect 5340 5496 5348 5504
rect 5388 5496 5396 5504
rect 5468 5496 5476 5504
rect 5628 5496 5636 5504
rect 5756 5496 5764 5504
rect 5852 5496 5860 5504
rect 5900 5496 5908 5504
rect 5996 5496 6004 5504
rect 6028 5496 6036 5504
rect 6188 5496 6196 5504
rect 6220 5496 6228 5504
rect 6252 5496 6260 5504
rect 6316 5496 6324 5504
rect 4732 5476 4740 5484
rect 4828 5476 4836 5484
rect 4892 5476 4900 5484
rect 4988 5476 4996 5484
rect 5116 5476 5124 5484
rect 5436 5476 5444 5484
rect 5548 5476 5556 5484
rect 5580 5476 5588 5484
rect 5756 5476 5764 5484
rect 5884 5476 5892 5484
rect 6044 5476 6052 5484
rect 6508 5496 6516 5504
rect 6540 5496 6548 5504
rect 6556 5496 6564 5504
rect 6620 5496 6628 5504
rect 6636 5496 6644 5504
rect 6684 5496 6692 5504
rect 6748 5496 6756 5504
rect 6828 5496 6836 5504
rect 6956 5496 6964 5504
rect 7132 5496 7140 5504
rect 7276 5496 7284 5504
rect 7420 5496 7428 5504
rect 7468 5496 7476 5504
rect 7692 5496 7700 5504
rect 7756 5494 7764 5502
rect 7868 5496 7876 5504
rect 7948 5496 7956 5504
rect 7996 5496 8004 5504
rect 8076 5496 8084 5504
rect 8108 5496 8116 5504
rect 6380 5476 6388 5484
rect 6476 5476 6484 5484
rect 6492 5476 6500 5484
rect 6572 5476 6580 5484
rect 6620 5476 6628 5484
rect 6636 5476 6644 5484
rect 6908 5476 6916 5484
rect 7260 5476 7268 5484
rect 7516 5476 7524 5484
rect 7964 5476 7972 5484
rect 7980 5476 7988 5484
rect 8124 5476 8132 5484
rect 316 5456 324 5464
rect 444 5456 452 5464
rect 604 5456 612 5464
rect 668 5456 676 5464
rect 940 5456 948 5464
rect 1164 5456 1172 5464
rect 1228 5456 1236 5464
rect 1484 5456 1492 5464
rect 1548 5456 1556 5464
rect 1804 5456 1812 5464
rect 1868 5456 1876 5464
rect 2028 5456 2036 5464
rect 2300 5456 2308 5464
rect 2316 5456 2324 5464
rect 2380 5456 2388 5464
rect 2764 5456 2772 5464
rect 3004 5456 3012 5464
rect 3516 5456 3524 5464
rect 4092 5456 4100 5464
rect 4124 5456 4132 5464
rect 4172 5456 4180 5464
rect 4204 5456 4212 5464
rect 4332 5456 4340 5464
rect 4748 5456 4756 5464
rect 5212 5456 5220 5464
rect 5500 5456 5508 5464
rect 5948 5456 5956 5464
rect 6108 5456 6116 5464
rect 6124 5456 6132 5464
rect 6188 5456 6196 5464
rect 6268 5456 6276 5464
rect 6700 5456 6708 5464
rect 6876 5456 6884 5464
rect 7084 5456 7092 5464
rect 7180 5456 7188 5464
rect 7244 5456 7252 5464
rect 7340 5456 7348 5464
rect 7548 5456 7556 5464
rect 7612 5456 7620 5464
rect 7820 5456 7828 5464
rect 8044 5456 8052 5464
rect 188 5436 196 5444
rect 236 5436 244 5444
rect 396 5436 404 5444
rect 684 5436 692 5444
rect 924 5436 932 5444
rect 1212 5436 1220 5444
rect 1756 5436 1764 5444
rect 1820 5436 1828 5444
rect 2060 5436 2068 5444
rect 2604 5436 2612 5444
rect 2828 5436 2836 5444
rect 2860 5436 2868 5444
rect 3132 5436 3140 5444
rect 3164 5436 3172 5444
rect 3420 5436 3428 5444
rect 3612 5436 3620 5444
rect 3836 5436 3844 5444
rect 3852 5436 3860 5444
rect 4236 5436 4244 5444
rect 4300 5436 4308 5444
rect 4412 5436 4420 5444
rect 5196 5436 5204 5444
rect 5276 5436 5284 5444
rect 5836 5436 5844 5444
rect 6284 5436 6292 5444
rect 6588 5436 6596 5444
rect 6796 5436 6804 5444
rect 7068 5436 7076 5444
rect 7100 5436 7108 5444
rect 7628 5436 7636 5444
rect 7836 5436 7844 5444
rect 8076 5436 8084 5444
rect 604 5416 612 5424
rect 1484 5416 1492 5424
rect 2316 5416 2324 5424
rect 6124 5416 6132 5424
rect 7244 5416 7252 5424
rect 7612 5416 7620 5424
rect 3278 5406 3286 5414
rect 3292 5406 3300 5414
rect 3306 5406 3314 5414
rect 6350 5406 6358 5414
rect 6364 5406 6372 5414
rect 6378 5406 6386 5414
rect 1596 5396 1604 5404
rect 4812 5396 4820 5404
rect 5964 5396 5972 5404
rect 12 5376 20 5384
rect 428 5376 436 5384
rect 796 5376 804 5384
rect 1132 5376 1140 5384
rect 1196 5376 1204 5384
rect 1404 5376 1412 5384
rect 1676 5376 1684 5384
rect 1836 5376 1844 5384
rect 1948 5376 1956 5384
rect 1980 5376 1988 5384
rect 2172 5376 2180 5384
rect 2828 5376 2836 5384
rect 3036 5376 3044 5384
rect 3100 5376 3108 5384
rect 3212 5376 3220 5384
rect 3628 5376 3636 5384
rect 3916 5376 3924 5384
rect 4620 5376 4628 5384
rect 4796 5376 4804 5384
rect 5004 5376 5012 5384
rect 5452 5376 5460 5384
rect 5708 5376 5716 5384
rect 6556 5376 6564 5384
rect 6636 5376 6644 5384
rect 6700 5376 6708 5384
rect 6764 5376 6772 5384
rect 7900 5376 7908 5384
rect 8012 5376 8020 5384
rect 204 5356 212 5364
rect 620 5356 628 5364
rect 636 5356 644 5364
rect 652 5356 660 5364
rect 1308 5356 1316 5364
rect 1596 5356 1604 5364
rect 1644 5356 1652 5364
rect 1692 5356 1700 5364
rect 1740 5356 1748 5364
rect 1964 5356 1972 5364
rect 1996 5356 2004 5364
rect 2028 5356 2036 5364
rect 2620 5356 2628 5364
rect 2636 5356 2644 5364
rect 3228 5356 3236 5364
rect 3516 5356 3524 5364
rect 4012 5356 4020 5364
rect 4028 5356 4036 5364
rect 4140 5356 4148 5364
rect 4284 5356 4292 5364
rect 4316 5356 4324 5364
rect 4812 5356 4820 5364
rect 4988 5356 4996 5364
rect 5180 5356 5188 5364
rect 5196 5356 5204 5364
rect 5292 5356 5300 5364
rect 5372 5356 5380 5364
rect 5516 5356 5524 5364
rect 5548 5356 5556 5364
rect 5900 5356 5908 5364
rect 5964 5356 5972 5364
rect 6316 5356 6324 5364
rect 6588 5356 6596 5364
rect 6620 5356 6628 5364
rect 6652 5356 6660 5364
rect 6780 5356 6788 5364
rect 7196 5356 7204 5364
rect 7324 5356 7332 5364
rect 7420 5356 7428 5364
rect 7484 5356 7492 5364
rect 7964 5356 7972 5364
rect 8028 5356 8036 5364
rect 124 5336 132 5344
rect 220 5336 228 5344
rect 284 5336 292 5344
rect 316 5336 324 5344
rect 348 5336 356 5344
rect 396 5336 404 5344
rect 412 5336 420 5344
rect 460 5336 468 5344
rect 476 5336 484 5344
rect 540 5336 548 5344
rect 620 5336 628 5344
rect 700 5336 708 5344
rect 716 5336 724 5344
rect 812 5336 820 5344
rect 844 5336 852 5344
rect 940 5336 948 5344
rect 972 5336 980 5344
rect 1148 5336 1156 5344
rect 1244 5336 1252 5344
rect 1292 5336 1300 5344
rect 1516 5336 1524 5344
rect 1900 5336 1908 5344
rect 2060 5336 2068 5344
rect 2092 5336 2100 5344
rect 2124 5336 2132 5344
rect 2204 5336 2212 5344
rect 2236 5336 2244 5344
rect 2268 5336 2276 5344
rect 2348 5336 2356 5344
rect 2412 5336 2420 5344
rect 2444 5336 2452 5344
rect 2668 5336 2676 5344
rect 2908 5336 2916 5344
rect 3084 5336 3092 5344
rect 3164 5336 3172 5344
rect 3324 5336 3332 5344
rect 3532 5336 3540 5344
rect 3548 5336 3556 5344
rect 3580 5336 3588 5344
rect 3644 5336 3652 5344
rect 3660 5336 3668 5344
rect 3692 5336 3700 5344
rect 4060 5336 4068 5344
rect 140 5318 148 5326
rect 252 5316 260 5324
rect 268 5316 276 5324
rect 300 5316 308 5324
rect 364 5316 372 5324
rect 460 5316 468 5324
rect 556 5316 564 5324
rect 828 5316 836 5324
rect 844 5316 852 5324
rect 1020 5316 1028 5324
rect 1356 5316 1364 5324
rect 1372 5316 1380 5324
rect 1500 5316 1508 5324
rect 1708 5316 1716 5324
rect 1916 5316 1924 5324
rect 2028 5316 2036 5324
rect 2076 5316 2084 5324
rect 2108 5316 2116 5324
rect 2140 5316 2148 5324
rect 2188 5316 2196 5324
rect 2220 5316 2228 5324
rect 2252 5316 2260 5324
rect 236 5296 244 5304
rect 316 5296 324 5304
rect 380 5296 388 5304
rect 428 5296 436 5304
rect 492 5296 500 5304
rect 524 5296 532 5304
rect 668 5296 676 5304
rect 764 5296 772 5304
rect 1260 5296 1268 5304
rect 1292 5296 1300 5304
rect 1388 5296 1396 5304
rect 2300 5296 2308 5304
rect 2332 5316 2340 5324
rect 2380 5316 2388 5324
rect 2396 5316 2404 5324
rect 2476 5318 2484 5326
rect 2700 5318 2708 5326
rect 2892 5318 2900 5326
rect 3068 5316 3076 5324
rect 3180 5316 3188 5324
rect 3356 5318 3364 5326
rect 3564 5316 3572 5324
rect 3676 5316 3684 5324
rect 3772 5318 3780 5326
rect 3820 5316 3828 5324
rect 3948 5316 3956 5324
rect 3980 5316 3988 5324
rect 4012 5316 4020 5324
rect 4108 5336 4116 5344
rect 4204 5336 4212 5344
rect 4220 5336 4228 5344
rect 4284 5336 4292 5344
rect 4332 5336 4340 5344
rect 4764 5336 4772 5344
rect 4924 5336 4932 5344
rect 5020 5336 5028 5344
rect 5116 5336 5124 5344
rect 5228 5336 5236 5344
rect 5244 5336 5252 5344
rect 5436 5336 5444 5344
rect 5500 5336 5508 5344
rect 5564 5336 5572 5344
rect 5996 5336 6004 5344
rect 6252 5336 6260 5344
rect 6380 5336 6388 5344
rect 6524 5336 6532 5344
rect 6572 5336 6580 5344
rect 6716 5336 6724 5344
rect 6796 5336 6804 5344
rect 7004 5336 7012 5344
rect 7068 5336 7076 5344
rect 7084 5336 7092 5344
rect 7132 5336 7140 5344
rect 7164 5336 7172 5344
rect 7244 5336 7252 5344
rect 7260 5336 7268 5344
rect 7356 5336 7364 5344
rect 7388 5336 7396 5344
rect 7516 5336 7524 5344
rect 7708 5336 7716 5344
rect 7740 5336 7748 5344
rect 7772 5336 7780 5344
rect 7868 5336 7876 5344
rect 7996 5336 8004 5344
rect 8028 5336 8036 5344
rect 8140 5336 8148 5344
rect 4092 5316 4100 5324
rect 4156 5316 4164 5324
rect 4188 5316 4196 5324
rect 4236 5316 4244 5324
rect 4252 5316 4260 5324
rect 4396 5316 4404 5324
rect 4428 5316 4436 5324
rect 4492 5318 4500 5326
rect 4556 5316 4564 5324
rect 4636 5316 4644 5324
rect 4780 5316 4788 5324
rect 4892 5316 4900 5324
rect 4908 5316 4916 5324
rect 4940 5316 4948 5324
rect 5068 5316 5076 5324
rect 5132 5316 5140 5324
rect 5148 5316 5156 5324
rect 5276 5316 5284 5324
rect 5340 5316 5348 5324
rect 5420 5316 5428 5324
rect 5484 5316 5492 5324
rect 5516 5316 5524 5324
rect 5692 5316 5700 5324
rect 5772 5316 5780 5324
rect 5836 5318 5844 5326
rect 6044 5316 6052 5324
rect 6076 5316 6084 5324
rect 6204 5316 6212 5324
rect 6268 5316 6276 5324
rect 6316 5316 6324 5324
rect 6444 5316 6452 5324
rect 6620 5316 6628 5324
rect 6732 5316 6740 5324
rect 6876 5316 6884 5324
rect 6924 5316 6932 5324
rect 7020 5316 7028 5324
rect 7116 5316 7124 5324
rect 7180 5316 7188 5324
rect 2364 5296 2372 5304
rect 3100 5296 3108 5304
rect 3212 5296 3220 5304
rect 3500 5296 3508 5304
rect 3596 5296 3604 5304
rect 3612 5296 3620 5304
rect 3708 5296 3716 5304
rect 3916 5296 3924 5304
rect 4268 5296 4276 5304
rect 4380 5296 4388 5304
rect 5052 5296 5060 5304
rect 5196 5296 5204 5304
rect 5948 5296 5956 5304
rect 6220 5296 6228 5304
rect 6332 5296 6340 5304
rect 6428 5296 6436 5304
rect 6492 5296 6500 5304
rect 6700 5296 6708 5304
rect 7020 5296 7028 5304
rect 7068 5296 7076 5304
rect 7100 5296 7108 5304
rect 7228 5316 7236 5324
rect 7292 5316 7300 5324
rect 7340 5316 7348 5324
rect 7404 5316 7412 5324
rect 7452 5316 7460 5324
rect 7564 5316 7572 5324
rect 7692 5316 7700 5324
rect 7756 5316 7764 5324
rect 7852 5316 7860 5324
rect 7900 5316 7908 5324
rect 7948 5316 7956 5324
rect 7980 5316 7988 5324
rect 8044 5316 8052 5324
rect 7772 5296 7780 5304
rect 7804 5296 7812 5304
rect 7884 5296 7892 5304
rect 556 5276 564 5284
rect 2604 5276 2612 5284
rect 2796 5276 2804 5284
rect 4876 5276 4884 5284
rect 6188 5276 6196 5284
rect 6460 5276 6468 5284
rect 6636 5276 6644 5284
rect 6988 5276 6996 5284
rect 7292 5276 7300 5284
rect 7820 5276 7828 5284
rect 7916 5276 7924 5284
rect 6172 5256 6180 5264
rect 7436 5256 7444 5264
rect 1612 5236 1620 5244
rect 3020 5236 3028 5244
rect 3244 5236 3252 5244
rect 3484 5236 3492 5244
rect 3900 5236 3908 5244
rect 3980 5236 3988 5244
rect 4140 5236 4148 5244
rect 5084 5236 5092 5244
rect 5148 5236 5156 5244
rect 5708 5236 5716 5244
rect 6156 5236 6164 5244
rect 6300 5236 6308 5244
rect 6444 5236 6452 5244
rect 7164 5236 7172 5244
rect 7388 5236 7396 5244
rect 7676 5236 7684 5244
rect 7740 5236 7748 5244
rect 7852 5236 7860 5244
rect 1742 5206 1750 5214
rect 1756 5206 1764 5214
rect 1770 5206 1778 5214
rect 4814 5206 4822 5214
rect 4828 5206 4836 5214
rect 4842 5206 4850 5214
rect 460 5176 468 5184
rect 908 5176 916 5184
rect 1804 5176 1812 5184
rect 4332 5176 4340 5184
rect 4380 5176 4388 5184
rect 4444 5176 4452 5184
rect 5292 5176 5300 5184
rect 5836 5176 5844 5184
rect 6140 5176 6148 5184
rect 6172 5176 6180 5184
rect 6540 5176 6548 5184
rect 7772 5176 7780 5184
rect 8012 5176 8020 5184
rect 4636 5156 4644 5164
rect 6236 5156 6244 5164
rect 6508 5156 6516 5164
rect 540 5136 548 5144
rect 668 5136 676 5144
rect 1308 5136 1316 5144
rect 1388 5136 1396 5144
rect 2028 5136 2036 5144
rect 2332 5136 2340 5144
rect 2540 5136 2548 5144
rect 2860 5136 2868 5144
rect 3212 5136 3220 5144
rect 3516 5136 3524 5144
rect 3788 5136 3796 5144
rect 4828 5136 4836 5144
rect 7116 5136 7124 5144
rect 7628 5136 7636 5144
rect 7884 5136 7892 5144
rect 1180 5116 1188 5124
rect 1276 5116 1284 5124
rect 1340 5116 1348 5124
rect 1356 5116 1364 5124
rect 76 5096 84 5104
rect 124 5096 132 5104
rect 204 5096 212 5104
rect 252 5096 260 5104
rect 268 5096 276 5104
rect 492 5096 500 5104
rect 604 5096 612 5104
rect 876 5096 884 5104
rect 988 5096 996 5104
rect 1116 5096 1124 5104
rect 1148 5096 1156 5104
rect 1212 5096 1220 5104
rect 1324 5096 1332 5104
rect 1372 5096 1380 5104
rect 1468 5094 1476 5102
rect 1516 5096 1524 5104
rect 1660 5094 1668 5102
rect 1916 5096 1924 5104
rect 2188 5116 2196 5124
rect 2252 5116 2260 5124
rect 2444 5116 2452 5124
rect 2556 5116 2564 5124
rect 2572 5116 2580 5124
rect 2588 5116 2596 5124
rect 2156 5096 2164 5104
rect 2236 5096 2244 5104
rect 2492 5096 2500 5104
rect 2620 5096 2628 5104
rect 2732 5094 2740 5102
rect 2796 5096 2804 5104
rect 2924 5116 2932 5124
rect 2956 5116 2964 5124
rect 3356 5116 3364 5124
rect 3004 5096 3012 5104
rect 3100 5096 3108 5104
rect 3260 5096 3268 5104
rect 3340 5096 3348 5104
rect 3420 5096 3428 5104
rect 3436 5096 3444 5104
rect 3468 5096 3476 5104
rect 3628 5116 3636 5124
rect 3724 5116 3732 5124
rect 3756 5116 3764 5124
rect 3852 5116 3860 5124
rect 3948 5116 3956 5124
rect 4732 5116 4740 5124
rect 4748 5116 4756 5124
rect 5004 5116 5012 5124
rect 5020 5116 5028 5124
rect 5404 5116 5412 5124
rect 5948 5116 5956 5124
rect 6204 5116 6212 5124
rect 6268 5116 6276 5124
rect 6412 5116 6420 5124
rect 6460 5116 6468 5124
rect 7068 5116 7076 5124
rect 3548 5096 3556 5104
rect 3580 5096 3588 5104
rect 3644 5096 3652 5104
rect 3660 5096 3668 5104
rect 3740 5096 3748 5104
rect 3788 5096 3796 5104
rect 3884 5096 3892 5104
rect 4012 5094 4020 5102
rect 4076 5096 4084 5104
rect 4204 5094 4212 5102
rect 4268 5096 4276 5104
rect 4524 5096 4532 5104
rect 4556 5096 4564 5104
rect 4700 5096 4708 5104
rect 4716 5096 4724 5104
rect 4876 5096 4884 5104
rect 4924 5096 4932 5104
rect 5036 5096 5044 5104
rect 5068 5096 5076 5104
rect 5164 5094 5172 5102
rect 5212 5096 5220 5104
rect 5388 5096 5396 5104
rect 5452 5096 5460 5104
rect 5596 5094 5604 5102
rect 5660 5096 5668 5104
rect 5788 5096 5796 5104
rect 5916 5096 5924 5104
rect 6028 5096 6036 5104
rect 6076 5096 6084 5104
rect 6172 5096 6180 5104
rect 6236 5096 6244 5104
rect 6284 5096 6292 5104
rect 6348 5096 6356 5104
rect 7132 5116 7140 5124
rect 7676 5116 7684 5124
rect 7708 5116 7716 5124
rect 7804 5116 7812 5124
rect 7996 5116 8004 5124
rect 8076 5116 8084 5124
rect 6700 5094 6708 5102
rect 6892 5094 6900 5102
rect 7164 5096 7172 5104
rect 7244 5096 7252 5104
rect 7292 5096 7300 5104
rect 7324 5096 7332 5104
rect 7340 5096 7348 5104
rect 7500 5096 7508 5104
rect 7676 5096 7684 5104
rect 7772 5096 7780 5104
rect 7852 5096 7860 5104
rect 7868 5096 7876 5104
rect 7932 5096 7940 5104
rect 7948 5096 7956 5104
rect 8044 5096 8052 5104
rect 8124 5096 8132 5104
rect 236 5076 244 5084
rect 268 5076 276 5084
rect 364 5076 372 5084
rect 572 5076 580 5084
rect 636 5076 644 5084
rect 684 5076 692 5084
rect 812 5076 820 5084
rect 1132 5076 1140 5084
rect 1228 5076 1236 5084
rect 1244 5076 1252 5084
rect 1308 5076 1316 5084
rect 1404 5076 1412 5084
rect 1628 5076 1636 5084
rect 1868 5076 1876 5084
rect 2140 5076 2148 5084
rect 2172 5076 2180 5084
rect 2220 5076 2228 5084
rect 2236 5076 2244 5084
rect 2300 5076 2308 5084
rect 2396 5076 2404 5084
rect 2476 5076 2484 5084
rect 2524 5076 2532 5084
rect 2540 5076 2548 5084
rect 2604 5076 2612 5084
rect 2876 5076 2884 5084
rect 2956 5076 2964 5084
rect 3020 5076 3028 5084
rect 3052 5076 3060 5084
rect 3372 5076 3380 5084
rect 3388 5080 3396 5088
rect 3452 5076 3460 5084
rect 3500 5076 3508 5084
rect 3516 5076 3524 5084
rect 3564 5076 3572 5084
rect 3676 5076 3684 5084
rect 3692 5076 3700 5084
rect 3724 5076 3732 5084
rect 3884 5076 3892 5084
rect 3900 5076 3908 5084
rect 3932 5076 3940 5084
rect 3980 5076 3988 5084
rect 4220 5076 4228 5084
rect 4476 5076 4484 5084
rect 4748 5076 4756 5084
rect 4780 5076 4788 5084
rect 4796 5076 4804 5084
rect 4908 5076 4916 5084
rect 4940 5076 4948 5084
rect 4972 5076 4980 5084
rect 5132 5076 5140 5084
rect 5260 5076 5268 5084
rect 204 5056 212 5064
rect 380 5056 388 5064
rect 444 5056 452 5064
rect 524 5056 532 5064
rect 556 5056 564 5064
rect 588 5056 596 5064
rect 972 5056 980 5064
rect 2044 5056 2052 5064
rect 2108 5056 2116 5064
rect 2188 5056 2196 5064
rect 2428 5056 2436 5064
rect 2444 5056 2452 5064
rect 2668 5056 2676 5064
rect 3228 5056 3236 5064
rect 3580 5056 3588 5064
rect 3612 5056 3620 5064
rect 3836 5056 3844 5064
rect 188 5036 196 5044
rect 396 5036 404 5044
rect 460 5036 468 5044
rect 508 5036 516 5044
rect 828 5036 836 5044
rect 1100 5036 1108 5044
rect 1260 5036 1268 5044
rect 1596 5036 1604 5044
rect 2092 5036 2100 5044
rect 2892 5036 2900 5044
rect 3868 5036 3876 5044
rect 4140 5036 4148 5044
rect 4332 5036 4340 5044
rect 4412 5056 4420 5064
rect 4652 5056 4660 5064
rect 5100 5056 5108 5064
rect 5308 5056 5316 5064
rect 5436 5076 5444 5084
rect 5564 5076 5572 5084
rect 5772 5076 5780 5084
rect 5932 5076 5940 5084
rect 6060 5076 6068 5084
rect 6156 5076 6164 5084
rect 6220 5076 6228 5084
rect 6300 5076 6308 5084
rect 6332 5076 6340 5084
rect 6460 5076 6468 5084
rect 6476 5076 6484 5084
rect 6492 5076 6500 5084
rect 6732 5076 6740 5084
rect 6828 5076 6836 5084
rect 6924 5076 6932 5084
rect 7036 5076 7044 5084
rect 7116 5076 7124 5084
rect 7228 5076 7236 5084
rect 7516 5076 7524 5084
rect 7916 5076 7924 5084
rect 7932 5076 7940 5084
rect 8028 5076 8036 5084
rect 8060 5076 8068 5084
rect 8092 5076 8100 5084
rect 4876 5036 4884 5044
rect 5356 5036 5364 5044
rect 5532 5056 5540 5064
rect 5756 5056 5764 5064
rect 5868 5056 5876 5064
rect 6316 5056 6324 5064
rect 6524 5056 6532 5064
rect 6556 5056 6564 5064
rect 6956 5056 6964 5064
rect 7020 5056 7028 5064
rect 7212 5056 7220 5064
rect 7356 5056 7364 5064
rect 7388 5056 7396 5064
rect 7420 5056 7428 5064
rect 7628 5056 7636 5064
rect 7724 5056 7732 5064
rect 7820 5056 7828 5064
rect 7996 5056 8004 5064
rect 5516 5036 5524 5044
rect 5740 5036 5748 5044
rect 5836 5036 5844 5044
rect 6412 5036 6420 5044
rect 6572 5036 6580 5044
rect 6764 5036 6772 5044
rect 7004 5036 7012 5044
rect 7132 5036 7140 5044
rect 7276 5036 7284 5044
rect 380 5016 388 5024
rect 2108 5016 2116 5024
rect 7020 5016 7028 5024
rect 7420 5016 7428 5024
rect 3278 5006 3286 5014
rect 3292 5006 3300 5014
rect 3306 5006 3314 5014
rect 6350 5006 6358 5014
rect 6364 5006 6372 5014
rect 6378 5006 6386 5014
rect 972 4976 980 4984
rect 1068 4976 1076 4984
rect 1116 4976 1124 4984
rect 1212 4976 1220 4984
rect 1372 4976 1380 4984
rect 2124 4976 2132 4984
rect 2732 4976 2740 4984
rect 3100 4976 3108 4984
rect 3260 4976 3268 4984
rect 3436 4976 3444 4984
rect 3612 4976 3620 4984
rect 3804 4976 3812 4984
rect 4636 4976 4644 4984
rect 4700 4976 4708 4984
rect 5228 4976 5236 4984
rect 5516 4976 5524 4984
rect 5548 4976 5556 4984
rect 5996 4976 6004 4984
rect 6764 4976 6772 4984
rect 6988 4976 6996 4984
rect 7052 4976 7060 4984
rect 7372 4976 7380 4984
rect 7420 4976 7428 4984
rect 7948 4976 7956 4984
rect 8076 4976 8084 4984
rect 12 4956 20 4964
rect 28 4956 36 4964
rect 460 4956 468 4964
rect 1180 4956 1188 4964
rect 1452 4956 1460 4964
rect 1484 4956 1492 4964
rect 1580 4956 1588 4964
rect 2220 4956 2228 4964
rect 2572 4956 2580 4964
rect 2668 4956 2676 4964
rect 2908 4956 2916 4964
rect 3116 4956 3124 4964
rect 3228 4956 3236 4964
rect 3388 4956 3396 4964
rect 3580 4956 3588 4964
rect 3740 4956 3748 4964
rect 3884 4956 3892 4964
rect 3900 4956 3908 4964
rect 3980 4956 3988 4964
rect 4124 4956 4132 4964
rect 4220 4956 4228 4964
rect 4444 4956 4452 4964
rect 4716 4956 4724 4964
rect 5132 4956 5140 4964
rect 44 4936 52 4944
rect 92 4936 100 4944
rect 124 4936 132 4944
rect 204 4936 212 4944
rect 268 4936 276 4944
rect 284 4936 292 4944
rect 412 4936 420 4944
rect 556 4936 564 4944
rect 652 4936 660 4944
rect 684 4936 692 4944
rect 860 4936 868 4944
rect 1004 4936 1012 4944
rect 1196 4936 1204 4944
rect 1228 4936 1236 4944
rect 1308 4936 1316 4944
rect 1420 4936 1428 4944
rect 1516 4936 1524 4944
rect 1548 4936 1556 4944
rect 1612 4936 1620 4944
rect 1804 4936 1812 4944
rect 1932 4936 1940 4944
rect 1964 4936 1972 4944
rect 2284 4936 2292 4944
rect 2300 4936 2308 4944
rect 2348 4936 2356 4944
rect 2428 4936 2436 4944
rect 2476 4936 2484 4944
rect 2524 4936 2532 4944
rect 2636 4936 2644 4944
rect 2684 4936 2692 4944
rect 2764 4936 2772 4944
rect 2796 4936 2804 4944
rect 3004 4936 3012 4944
rect 3228 4936 3236 4944
rect 3276 4936 3284 4944
rect 3420 4936 3428 4944
rect 3500 4936 3508 4944
rect 4588 4936 4596 4944
rect 4668 4932 4676 4940
rect 4748 4936 4756 4944
rect 4972 4936 4980 4944
rect 5068 4936 5076 4944
rect 5404 4936 5412 4944
rect 5532 4936 5540 4944
rect 5868 4956 5876 4964
rect 6636 4956 6644 4964
rect 6812 4956 6820 4964
rect 7004 4956 7012 4964
rect 7388 4956 7396 4964
rect 7740 4956 7748 4964
rect 8108 4956 8116 4964
rect 5644 4936 5652 4944
rect 5740 4936 5748 4944
rect 5964 4936 5972 4944
rect 6028 4936 6036 4944
rect 6060 4936 6068 4944
rect 6300 4936 6308 4944
rect 6332 4936 6340 4944
rect 6428 4936 6436 4944
rect 6668 4936 6676 4944
rect 6748 4936 6756 4944
rect 6780 4936 6788 4944
rect 6844 4936 6852 4944
rect 6860 4936 6868 4944
rect 6924 4936 6932 4944
rect 6972 4936 6980 4944
rect 7084 4936 7092 4944
rect 7180 4936 7188 4944
rect 7260 4936 7268 4944
rect 7516 4936 7524 4944
rect 7676 4936 7684 4944
rect 7820 4936 7828 4944
rect 7884 4936 7892 4944
rect 7932 4936 7940 4944
rect 7980 4932 7988 4940
rect 7996 4936 8004 4944
rect 8012 4936 8020 4944
rect 8092 4936 8100 4944
rect 172 4916 180 4924
rect 188 4916 196 4924
rect 268 4916 276 4924
rect 364 4916 372 4924
rect 412 4916 420 4924
rect 508 4916 516 4924
rect 556 4916 564 4924
rect 604 4916 612 4924
rect 636 4916 644 4924
rect 716 4918 724 4926
rect 1148 4916 1156 4924
rect 1196 4916 1204 4924
rect 1260 4916 1268 4924
rect 1324 4916 1332 4924
rect 76 4896 84 4904
rect 140 4896 148 4904
rect 156 4896 164 4904
rect 220 4896 228 4904
rect 252 4896 260 4904
rect 316 4896 324 4904
rect 380 4896 388 4904
rect 396 4896 404 4904
rect 588 4896 596 4904
rect 604 4896 612 4904
rect 636 4896 644 4904
rect 1228 4896 1236 4904
rect 1356 4896 1364 4904
rect 1500 4916 1508 4924
rect 2012 4916 2020 4924
rect 2156 4916 2164 4924
rect 2252 4916 2260 4924
rect 2268 4916 2276 4924
rect 2332 4916 2340 4924
rect 2380 4916 2388 4924
rect 2444 4916 2452 4924
rect 2476 4916 2484 4924
rect 2572 4916 2580 4924
rect 2588 4916 2596 4924
rect 2636 4916 2644 4924
rect 2700 4916 2708 4924
rect 2748 4916 2756 4924
rect 2780 4916 2788 4924
rect 2812 4916 2820 4924
rect 2876 4916 2884 4924
rect 2972 4918 2980 4926
rect 3148 4916 3156 4924
rect 3180 4916 3188 4924
rect 3356 4916 3364 4924
rect 1436 4896 1444 4904
rect 2140 4896 2148 4904
rect 2220 4896 2228 4904
rect 2236 4896 2244 4904
rect 2300 4896 2308 4904
rect 2364 4896 2372 4904
rect 2460 4896 2468 4904
rect 2652 4896 2660 4904
rect 2828 4896 2836 4904
rect 2860 4896 2868 4904
rect 3148 4896 3156 4904
rect 3292 4896 3300 4904
rect 3340 4896 3348 4904
rect 3388 4896 3396 4904
rect 3548 4916 3556 4924
rect 3740 4918 3748 4926
rect 3852 4916 3860 4924
rect 3980 4918 3988 4926
rect 4156 4916 4164 4924
rect 4252 4916 4260 4924
rect 4364 4916 4372 4924
rect 4412 4916 4420 4924
rect 4604 4916 4612 4924
rect 4940 4918 4948 4926
rect 5132 4918 5140 4926
rect 5196 4916 5204 4924
rect 5372 4918 5380 4926
rect 5452 4916 5460 4924
rect 5580 4916 5588 4924
rect 5756 4916 5764 4924
rect 5932 4918 5940 4926
rect 6108 4916 6116 4924
rect 6284 4916 6292 4924
rect 6396 4916 6404 4924
rect 6492 4918 6500 4926
rect 6540 4916 6548 4924
rect 6668 4916 6676 4924
rect 6700 4916 6708 4924
rect 6732 4916 6740 4924
rect 6796 4916 6804 4924
rect 6924 4916 6932 4924
rect 6956 4916 6964 4924
rect 7036 4916 7044 4924
rect 7116 4916 7124 4924
rect 7244 4918 7252 4926
rect 7548 4918 7556 4926
rect 7628 4916 7636 4924
rect 7660 4916 7668 4924
rect 7676 4916 7684 4924
rect 7772 4916 7780 4924
rect 7804 4916 7812 4924
rect 3468 4896 3476 4904
rect 3564 4896 3572 4904
rect 3804 4896 3812 4904
rect 4364 4896 4372 4904
rect 5436 4896 5444 4904
rect 5548 4896 5556 4904
rect 5692 4896 5700 4904
rect 5724 4896 5732 4904
rect 5756 4896 5764 4904
rect 6316 4896 6324 4904
rect 6428 4896 6436 4904
rect 6588 4896 6596 4904
rect 6876 4896 6884 4904
rect 6924 4896 6932 4904
rect 7020 4896 7028 4904
rect 7612 4896 7620 4904
rect 7692 4896 7700 4904
rect 7724 4896 7732 4904
rect 7772 4896 7780 4904
rect 7836 4896 7844 4904
rect 7900 4896 7908 4904
rect 8044 4896 8052 4904
rect 348 4876 356 4884
rect 428 4876 436 4884
rect 556 4876 564 4884
rect 1292 4876 1300 4884
rect 2092 4876 2100 4884
rect 2140 4876 2148 4884
rect 300 4856 308 4864
rect 844 4856 852 4864
rect 1468 4856 1476 4864
rect 2172 4876 2180 4884
rect 2396 4876 2404 4884
rect 2524 4876 2532 4884
rect 3420 4876 3428 4884
rect 3532 4876 3540 4884
rect 4716 4876 4724 4884
rect 4796 4876 4804 4884
rect 5468 4876 5476 4884
rect 5500 4876 5508 4884
rect 5996 4876 6004 4884
rect 6220 4876 6228 4884
rect 6620 4876 6628 4884
rect 6668 4876 6676 4884
rect 6908 4876 6916 4884
rect 7052 4876 7060 4884
rect 7644 4876 7652 4884
rect 8092 4876 8100 4884
rect 2380 4856 2388 4864
rect 5452 4856 5460 4864
rect 364 4836 372 4844
rect 476 4836 484 4844
rect 972 4836 980 4844
rect 1260 4836 1268 4844
rect 1548 4836 1556 4844
rect 1596 4836 1604 4844
rect 1724 4836 1732 4844
rect 3132 4836 3140 4844
rect 3548 4836 3556 4844
rect 3596 4836 3604 4844
rect 3916 4836 3924 4844
rect 4108 4836 4116 4844
rect 4156 4836 4164 4844
rect 4348 4836 4356 4844
rect 4476 4836 4484 4844
rect 5004 4836 5012 4844
rect 5244 4836 5252 4844
rect 5708 4836 5716 4844
rect 7404 4836 7412 4844
rect 7868 4836 7876 4844
rect 1742 4806 1750 4814
rect 1756 4806 1764 4814
rect 1770 4806 1778 4814
rect 4814 4806 4822 4814
rect 4828 4806 4836 4814
rect 4842 4806 4850 4814
rect 380 4776 388 4784
rect 892 4776 900 4784
rect 1196 4776 1204 4784
rect 3132 4776 3140 4784
rect 3292 4776 3300 4784
rect 3740 4776 3748 4784
rect 3884 4776 3892 4784
rect 4428 4776 4436 4784
rect 5148 4776 5156 4784
rect 5372 4776 5380 4784
rect 5548 4776 5556 4784
rect 5676 4776 5684 4784
rect 5820 4776 5828 4784
rect 6332 4776 6340 4784
rect 6572 4776 6580 4784
rect 6988 4776 6996 4784
rect 7692 4776 7700 4784
rect 764 4756 772 4764
rect 2860 4756 2868 4764
rect 5116 4756 5124 4764
rect 6892 4756 6900 4764
rect 588 4736 596 4744
rect 668 4736 676 4744
rect 1820 4736 1828 4744
rect 2124 4736 2132 4744
rect 2588 4736 2596 4744
rect 2828 4736 2836 4744
rect 3724 4736 3732 4744
rect 3772 4736 3780 4744
rect 4348 4736 4356 4744
rect 4636 4736 4644 4744
rect 4972 4736 4980 4744
rect 5164 4736 5172 4744
rect 5276 4736 5284 4744
rect 5692 4736 5700 4744
rect 5964 4736 5972 4744
rect 6076 4736 6084 4744
rect 6732 4736 6740 4744
rect 7404 4736 7412 4744
rect 7708 4736 7716 4744
rect 7884 4736 7892 4744
rect 284 4716 292 4724
rect 604 4716 612 4724
rect 652 4716 660 4724
rect 684 4716 692 4724
rect 1388 4716 1396 4724
rect 1452 4716 1460 4724
rect 140 4694 148 4702
rect 252 4696 260 4704
rect 268 4696 276 4704
rect 300 4696 308 4704
rect 364 4696 372 4704
rect 460 4694 468 4702
rect 524 4696 532 4704
rect 700 4696 708 4704
rect 748 4696 756 4704
rect 812 4696 820 4704
rect 828 4696 836 4704
rect 972 4694 980 4702
rect 1260 4696 1268 4704
rect 1548 4716 1556 4724
rect 1900 4716 1908 4724
rect 2156 4716 2164 4724
rect 2172 4716 2180 4724
rect 2796 4716 2804 4724
rect 3052 4716 3060 4724
rect 3580 4716 3588 4724
rect 3644 4716 3652 4724
rect 3692 4716 3700 4724
rect 1324 4694 1332 4702
rect 1596 4696 1604 4704
rect 1644 4696 1652 4704
rect 1708 4696 1716 4704
rect 172 4676 180 4684
rect 316 4676 324 4684
rect 348 4676 356 4684
rect 636 4676 644 4684
rect 652 4676 660 4684
rect 812 4676 820 4684
rect 860 4680 868 4688
rect 876 4676 884 4684
rect 940 4676 948 4684
rect 1308 4676 1316 4684
rect 1436 4676 1444 4684
rect 1484 4676 1492 4684
rect 1500 4676 1508 4684
rect 1580 4676 1588 4684
rect 1980 4696 1988 4704
rect 2044 4694 2052 4702
rect 2108 4696 2116 4704
rect 2284 4696 2292 4704
rect 2364 4696 2372 4704
rect 2380 4696 2388 4704
rect 2412 4696 2420 4704
rect 2444 4696 2452 4704
rect 2524 4696 2532 4704
rect 2588 4696 2596 4704
rect 2668 4696 2676 4704
rect 2732 4694 2740 4702
rect 2828 4696 2836 4704
rect 2924 4696 2932 4704
rect 2972 4696 2980 4704
rect 3116 4696 3124 4704
rect 3164 4696 3172 4704
rect 3196 4696 3204 4704
rect 3356 4696 3364 4704
rect 3420 4694 3428 4702
rect 3484 4696 3492 4704
rect 3516 4696 3524 4704
rect 3708 4696 3716 4704
rect 3772 4696 3780 4704
rect 3820 4716 3828 4724
rect 3932 4716 3940 4724
rect 4156 4716 4164 4724
rect 4444 4716 4452 4724
rect 3996 4696 4004 4704
rect 4012 4696 4020 4704
rect 4220 4694 4228 4702
rect 4284 4696 4292 4704
rect 4396 4696 4404 4704
rect 4476 4696 4484 4704
rect 4556 4696 4564 4704
rect 4860 4716 4868 4724
rect 4940 4716 4948 4724
rect 5004 4716 5012 4724
rect 5068 4716 5076 4724
rect 4668 4696 4676 4704
rect 4684 4696 4692 4704
rect 4732 4696 4740 4704
rect 4748 4696 4756 4704
rect 4828 4696 4836 4704
rect 4988 4696 4996 4704
rect 1804 4680 1812 4688
rect 1820 4676 1828 4684
rect 1852 4676 1860 4684
rect 2108 4676 2116 4684
rect 2220 4676 2228 4684
rect 2236 4676 2244 4684
rect 2396 4676 2404 4684
rect 2428 4676 2436 4684
rect 2524 4676 2532 4684
rect 2540 4676 2548 4684
rect 2764 4676 2772 4684
rect 2844 4676 2852 4684
rect 3020 4676 3028 4684
rect 3180 4676 3188 4684
rect 3228 4676 3236 4684
rect 3500 4676 3508 4684
rect 3564 4676 3572 4684
rect 3628 4676 3636 4684
rect 3676 4676 3684 4684
rect 3756 4676 3764 4684
rect 3868 4676 3876 4684
rect 3964 4676 3972 4684
rect 3980 4676 3988 4684
rect 4012 4676 4020 4684
rect 4108 4676 4116 4684
rect 4124 4676 4132 4684
rect 4364 4676 4372 4684
rect 4412 4676 4420 4684
rect 4460 4676 4468 4684
rect 4556 4676 4564 4684
rect 4572 4676 4580 4684
rect 4604 4676 4612 4684
rect 4620 4676 4628 4684
rect 4684 4676 4692 4684
rect 4764 4676 4772 4684
rect 4908 4676 4916 4684
rect 4988 4676 4996 4684
rect 5036 4696 5044 4704
rect 5196 4716 5204 4724
rect 5388 4716 5396 4724
rect 5484 4716 5492 4724
rect 5116 4696 5124 4704
rect 5180 4696 5188 4704
rect 5324 4696 5332 4704
rect 5516 4696 5524 4704
rect 5548 4696 5556 4704
rect 5596 4716 5604 4724
rect 5660 4716 5668 4724
rect 5756 4716 5764 4724
rect 5932 4716 5940 4724
rect 6092 4716 6100 4724
rect 6412 4716 6420 4724
rect 5628 4696 5636 4704
rect 5676 4696 5684 4704
rect 5772 4696 5780 4704
rect 5852 4696 5860 4704
rect 5932 4696 5940 4704
rect 6012 4696 6020 4704
rect 6028 4696 6036 4704
rect 6044 4696 6052 4704
rect 6156 4696 6164 4704
rect 6172 4696 6180 4704
rect 6236 4696 6244 4704
rect 6316 4696 6324 4704
rect 6524 4696 6532 4704
rect 6588 4696 6596 4704
rect 6652 4716 6660 4724
rect 6860 4716 6868 4724
rect 6956 4716 6964 4724
rect 7020 4716 7028 4724
rect 7036 4716 7044 4724
rect 6700 4696 6708 4704
rect 6748 4696 6756 4704
rect 6796 4696 6804 4704
rect 6924 4696 6932 4704
rect 6956 4696 6964 4704
rect 6988 4696 6996 4704
rect 7052 4696 7060 4704
rect 7068 4696 7076 4704
rect 7436 4716 7444 4724
rect 7292 4696 7300 4704
rect 7436 4696 7444 4704
rect 7484 4716 7492 4724
rect 7692 4716 7700 4724
rect 7852 4716 7860 4724
rect 8060 4716 8068 4724
rect 7516 4696 7524 4704
rect 7548 4696 7556 4704
rect 7628 4696 7636 4704
rect 7660 4696 7668 4704
rect 7692 4696 7700 4704
rect 7740 4696 7748 4704
rect 7804 4696 7812 4704
rect 7948 4696 7956 4704
rect 8012 4696 8020 4704
rect 5132 4676 5140 4684
rect 5212 4676 5220 4684
rect 5324 4676 5332 4684
rect 5340 4676 5348 4684
rect 5436 4676 5444 4684
rect 5452 4676 5460 4684
rect 5532 4676 5540 4684
rect 5644 4676 5652 4684
rect 5724 4676 5732 4684
rect 5740 4676 5748 4684
rect 5788 4676 5796 4684
rect 5820 4676 5828 4684
rect 6140 4676 6148 4684
rect 6220 4676 6228 4684
rect 6284 4676 6292 4684
rect 6444 4676 6452 4684
rect 6460 4676 6468 4684
rect 6476 4680 6484 4688
rect 6540 4676 6548 4684
rect 6572 4676 6580 4684
rect 6604 4676 6612 4684
rect 6684 4676 6692 4684
rect 6908 4676 6916 4684
rect 6972 4676 6980 4684
rect 7084 4676 7092 4684
rect 7132 4676 7140 4684
rect 7244 4676 7252 4684
rect 7420 4676 7428 4684
rect 7532 4676 7540 4684
rect 7564 4676 7572 4684
rect 7596 4676 7604 4684
rect 7612 4676 7620 4684
rect 7756 4676 7764 4684
rect 7788 4676 7796 4684
rect 7884 4676 7892 4684
rect 7996 4676 8004 4684
rect 8028 4676 8036 4684
rect 8124 4676 8132 4684
rect 204 4656 212 4664
rect 316 4656 324 4664
rect 396 4656 404 4664
rect 732 4656 740 4664
rect 908 4656 916 4664
rect 1116 4656 1124 4664
rect 1180 4656 1188 4664
rect 1388 4656 1396 4664
rect 1532 4656 1540 4664
rect 1628 4656 1636 4664
rect 1852 4656 1860 4664
rect 2252 4656 2260 4664
rect 2300 4656 2308 4664
rect 2364 4656 2372 4664
rect 2460 4656 2468 4664
rect 2492 4656 2500 4664
rect 3068 4656 3076 4664
rect 3532 4656 3540 4664
rect 3548 4656 3556 4664
rect 3580 4656 3588 4664
rect 3900 4656 3908 4664
rect 3916 4656 3924 4664
rect 3948 4656 3956 4664
rect 4524 4656 4532 4664
rect 4700 4656 4708 4664
rect 4924 4656 4932 4664
rect 5500 4656 5508 4664
rect 5884 4656 5892 4664
rect 6140 4656 6148 4664
rect 6204 4656 6212 4664
rect 6396 4656 6404 4664
rect 6796 4656 6804 4664
rect 6828 4656 6836 4664
rect 6876 4656 6884 4664
rect 7100 4656 7108 4664
rect 7148 4656 7156 4664
rect 7212 4656 7220 4664
rect 7628 4656 7636 4664
rect 7836 4656 7844 4664
rect 7852 4656 7860 4664
rect 7916 4656 7924 4664
rect 7948 4656 7956 4664
rect 7964 4656 7972 4664
rect 12 4636 20 4644
rect 1100 4636 1108 4644
rect 1164 4636 1172 4644
rect 1676 4636 1684 4644
rect 1900 4636 1908 4644
rect 1916 4636 1924 4644
rect 2476 4636 2484 4644
rect 2860 4636 2868 4644
rect 3084 4636 3092 4644
rect 4156 4636 4164 4644
rect 4508 4636 4516 4644
rect 4588 4636 4596 4644
rect 4780 4636 4788 4644
rect 5868 4636 5876 4644
rect 5916 4636 5924 4644
rect 6108 4636 6116 4644
rect 6188 4636 6196 4644
rect 6268 4636 6276 4644
rect 6364 4636 6372 4644
rect 6508 4636 6516 4644
rect 6620 4636 6628 4644
rect 6780 4636 6788 4644
rect 7196 4636 7204 4644
rect 7564 4636 7572 4644
rect 7772 4636 7780 4644
rect 7980 4636 7988 4644
rect 1180 4616 1188 4624
rect 7212 4616 7220 4624
rect 3278 4606 3286 4614
rect 3292 4606 3300 4614
rect 3306 4606 3314 4614
rect 6350 4606 6358 4614
rect 6364 4606 6372 4614
rect 6378 4606 6386 4614
rect 3420 4596 3428 4604
rect 3580 4596 3588 4604
rect 5244 4596 5252 4604
rect 252 4576 260 4584
rect 812 4576 820 4584
rect 860 4576 868 4584
rect 1324 4576 1332 4584
rect 2076 4576 2084 4584
rect 2124 4576 2132 4584
rect 2140 4576 2148 4584
rect 2780 4576 2788 4584
rect 2828 4576 2836 4584
rect 3228 4576 3236 4584
rect 3292 4576 3300 4584
rect 3500 4576 3508 4584
rect 3596 4576 3604 4584
rect 3692 4576 3700 4584
rect 3916 4576 3924 4584
rect 4236 4576 4244 4584
rect 4508 4576 4516 4584
rect 4652 4576 4660 4584
rect 4748 4576 4756 4584
rect 5260 4576 5268 4584
rect 5500 4576 5508 4584
rect 5708 4576 5716 4584
rect 5788 4576 5796 4584
rect 5932 4576 5940 4584
rect 7356 4576 7364 4584
rect 7564 4576 7572 4584
rect 7948 4576 7956 4584
rect 300 4556 308 4564
rect 348 4556 356 4564
rect 620 4556 628 4564
rect 956 4556 964 4564
rect 1004 4556 1012 4564
rect 1132 4556 1140 4564
rect 1596 4556 1604 4564
rect 1612 4556 1620 4564
rect 1740 4556 1748 4564
rect 172 4536 180 4544
rect 2060 4556 2068 4564
rect 2588 4556 2596 4564
rect 2748 4556 2756 4564
rect 2764 4556 2772 4564
rect 3036 4556 3044 4564
rect 3324 4556 3332 4564
rect 3420 4556 3428 4564
rect 3564 4556 3572 4564
rect 3580 4556 3588 4564
rect 3820 4556 3828 4564
rect 3852 4556 3860 4564
rect 4108 4556 4116 4564
rect 4220 4556 4228 4564
rect 4316 4556 4324 4564
rect 4732 4556 4740 4564
rect 4764 4556 4772 4564
rect 5084 4556 5092 4564
rect 5100 4556 5108 4564
rect 5228 4556 5236 4564
rect 5244 4556 5252 4564
rect 5308 4556 5316 4564
rect 5692 4556 5700 4564
rect 5724 4556 5732 4564
rect 6620 4556 6628 4564
rect 6636 4556 6644 4564
rect 6748 4556 6756 4564
rect 6780 4556 6788 4564
rect 6828 4556 6836 4564
rect 7164 4556 7172 4564
rect 412 4536 420 4544
rect 428 4536 436 4544
rect 508 4536 516 4544
rect 716 4536 724 4544
rect 844 4536 852 4544
rect 1292 4532 1300 4540
rect 1500 4536 1508 4544
rect 1532 4536 1540 4544
rect 1580 4536 1588 4544
rect 1612 4536 1620 4544
rect 1980 4536 1988 4544
rect 2092 4536 2100 4544
rect 2300 4536 2308 4544
rect 2396 4536 2404 4544
rect 2524 4536 2532 4544
rect 2716 4536 2724 4544
rect 2796 4536 2804 4544
rect 2860 4536 2868 4544
rect 2876 4536 2884 4544
rect 2972 4536 2980 4544
rect 3180 4536 3188 4544
rect 3244 4536 3252 4544
rect 3420 4536 3428 4544
rect 3532 4536 3540 4544
rect 3740 4536 3748 4544
rect 3772 4536 3780 4544
rect 3820 4536 3828 4544
rect 3900 4536 3908 4544
rect 3948 4536 3956 4544
rect 4028 4536 4036 4544
rect 4092 4536 4100 4544
rect 4172 4536 4180 4544
rect 4348 4536 4356 4544
rect 4524 4536 4532 4544
rect 4620 4536 4628 4544
rect 4636 4536 4644 4544
rect 4716 4536 4724 4544
rect 5004 4536 5012 4544
rect 5052 4536 5060 4544
rect 5116 4536 5124 4544
rect 5132 4536 5140 4544
rect 5180 4536 5188 4544
rect 5516 4536 5524 4544
rect 5548 4536 5556 4544
rect 5612 4536 5620 4544
rect 5756 4536 5764 4544
rect 5772 4536 5780 4544
rect 5804 4536 5812 4544
rect 5884 4536 5892 4544
rect 6044 4536 6052 4544
rect 6156 4536 6164 4544
rect 6172 4536 6180 4544
rect 6252 4536 6260 4544
rect 6492 4536 6500 4544
rect 6524 4536 6532 4544
rect 6540 4536 6548 4544
rect 6604 4536 6612 4544
rect 6764 4536 6772 4544
rect 6812 4536 6820 4544
rect 6908 4536 6916 4544
rect 6940 4536 6948 4544
rect 7132 4536 7140 4544
rect 7196 4536 7204 4544
rect 7244 4536 7252 4544
rect 7372 4536 7380 4544
rect 7420 4536 7428 4544
rect 7468 4536 7476 4544
rect 7484 4536 7492 4544
rect 7548 4536 7556 4544
rect 7580 4536 7588 4544
rect 7644 4536 7652 4544
rect 7676 4536 7684 4544
rect 7708 4536 7716 4544
rect 7740 4536 7748 4544
rect 7916 4536 7924 4544
rect 92 4516 100 4524
rect 204 4516 212 4524
rect 220 4516 228 4524
rect 300 4516 308 4524
rect 364 4516 372 4524
rect 380 4516 388 4524
rect 444 4516 452 4524
rect 524 4516 532 4524
rect 556 4516 564 4524
rect 684 4518 692 4526
rect 828 4516 836 4524
rect 940 4516 948 4524
rect 988 4516 996 4524
rect 1036 4516 1044 4524
rect 1068 4516 1076 4524
rect 1132 4518 1140 4526
rect 1276 4516 1284 4524
rect 1468 4518 1476 4526
rect 1548 4516 1556 4524
rect 1692 4516 1700 4524
rect 1740 4516 1748 4524
rect 1996 4518 2004 4526
rect 2204 4516 2212 4524
rect 2268 4518 2276 4526
rect 2332 4516 2340 4524
rect 2364 4516 2372 4524
rect 2412 4516 2420 4524
rect 2492 4516 2500 4524
rect 2540 4516 2548 4524
rect 2636 4516 2644 4524
rect 2652 4516 2660 4524
rect 2668 4516 2676 4524
rect 2812 4516 2820 4524
rect 3036 4518 3044 4526
rect 3196 4516 3204 4524
rect 3260 4516 3268 4524
rect 3580 4516 3588 4524
rect 3612 4516 3620 4524
rect 3660 4516 3668 4524
rect 3724 4516 3732 4524
rect 3788 4516 3796 4524
rect 3916 4516 3924 4524
rect 3980 4516 3988 4524
rect 4028 4516 4036 4524
rect 4124 4516 4132 4524
rect 4188 4516 4196 4524
rect 4268 4516 4276 4524
rect 4380 4518 4388 4526
rect 4972 4518 4980 4526
rect 316 4496 324 4504
rect 412 4496 420 4504
rect 476 4496 484 4504
rect 540 4496 548 4504
rect 892 4496 900 4504
rect 1020 4496 1028 4504
rect 1580 4496 1588 4504
rect 2124 4496 2132 4504
rect 2380 4496 2388 4504
rect 2444 4496 2452 4504
rect 2460 4496 2468 4504
rect 2508 4496 2516 4504
rect 2668 4496 2676 4504
rect 2684 4496 2692 4504
rect 2716 4496 2724 4504
rect 2828 4496 2836 4504
rect 3228 4496 3236 4504
rect 3308 4496 3316 4504
rect 3404 4496 3412 4504
rect 3676 4496 3684 4504
rect 3756 4496 3764 4504
rect 3852 4496 3860 4504
rect 3916 4496 3924 4504
rect 3964 4496 3972 4504
rect 4172 4496 4180 4504
rect 4220 4496 4228 4504
rect 4556 4496 4564 4504
rect 5036 4516 5044 4524
rect 5068 4516 5076 4524
rect 4684 4496 4692 4504
rect 5164 4496 5172 4504
rect 5388 4516 5396 4524
rect 5420 4516 5428 4524
rect 5532 4516 5540 4524
rect 5564 4516 5572 4524
rect 5612 4516 5620 4524
rect 5676 4516 5684 4524
rect 5756 4516 5764 4524
rect 5820 4516 5828 4524
rect 5836 4516 5844 4524
rect 5884 4516 5892 4524
rect 6060 4518 6068 4526
rect 6204 4516 6212 4524
rect 6284 4518 6292 4526
rect 6476 4516 6484 4524
rect 6604 4516 6612 4524
rect 6652 4516 6660 4524
rect 6684 4516 6692 4524
rect 6700 4516 6708 4524
rect 6796 4516 6804 4524
rect 6860 4516 6868 4524
rect 6972 4518 6980 4526
rect 7116 4516 7124 4524
rect 7164 4516 7172 4524
rect 7228 4518 7236 4526
rect 7500 4516 7508 4524
rect 7532 4516 7540 4524
rect 5564 4496 5572 4504
rect 5580 4496 5588 4504
rect 5628 4496 5636 4504
rect 5916 4496 5924 4504
rect 6124 4496 6132 4504
rect 6220 4496 6228 4504
rect 6556 4496 6564 4504
rect 6668 4496 6676 4504
rect 6876 4496 6884 4504
rect 7372 4496 7380 4504
rect 7436 4496 7444 4504
rect 7580 4496 7588 4504
rect 7724 4516 7732 4524
rect 7852 4516 7860 4524
rect 8012 4516 8020 4524
rect 8060 4516 8068 4524
rect 7644 4496 7652 4504
rect 7692 4496 7700 4504
rect 300 4476 308 4484
rect 444 4476 452 4484
rect 508 4476 516 4484
rect 1052 4476 1060 4484
rect 1372 4476 1380 4484
rect 2348 4476 2356 4484
rect 2412 4476 2420 4484
rect 2476 4476 2484 4484
rect 2540 4476 2548 4484
rect 2908 4476 2916 4484
rect 3132 4476 3140 4484
rect 3644 4476 3652 4484
rect 3948 4476 3956 4484
rect 3996 4476 4004 4484
rect 4076 4476 4084 4484
rect 4876 4476 4884 4484
rect 6412 4476 6420 4484
rect 6524 4476 6532 4484
rect 7100 4476 7108 4484
rect 7788 4476 7796 4484
rect 12 4436 20 4444
rect 252 4436 260 4444
rect 588 4436 596 4444
rect 972 4436 980 4444
rect 1260 4436 1268 4444
rect 1340 4436 1348 4444
rect 1804 4436 1812 4444
rect 1836 4436 1844 4444
rect 3164 4436 3172 4444
rect 3660 4436 3668 4444
rect 3836 4436 3844 4444
rect 4044 4436 4052 4444
rect 4780 4436 4788 4444
rect 4844 4436 4852 4444
rect 5868 4436 5876 4444
rect 5932 4436 5940 4444
rect 7756 4436 7764 4444
rect 7948 4436 7956 4444
rect 1742 4406 1750 4414
rect 1756 4406 1764 4414
rect 1770 4406 1778 4414
rect 4814 4406 4822 4414
rect 4828 4406 4836 4414
rect 4842 4406 4850 4414
rect 396 4376 404 4384
rect 860 4376 868 4384
rect 1084 4376 1092 4384
rect 1132 4376 1140 4384
rect 1468 4376 1476 4384
rect 2044 4376 2052 4384
rect 2796 4376 2804 4384
rect 2924 4376 2932 4384
rect 3308 4376 3316 4384
rect 3436 4376 3444 4384
rect 3516 4376 3524 4384
rect 3740 4376 3748 4384
rect 4092 4376 4100 4384
rect 4300 4376 4308 4384
rect 4348 4376 4356 4384
rect 4460 4376 4468 4384
rect 5292 4376 5300 4384
rect 5324 4376 5332 4384
rect 6108 4376 6116 4384
rect 6476 4376 6484 4384
rect 6604 4376 6612 4384
rect 6636 4376 6644 4384
rect 8028 4376 8036 4384
rect 8044 4376 8052 4384
rect 3004 4356 3012 4364
rect 3948 4356 3956 4364
rect 5580 4356 5588 4364
rect 7628 4356 7636 4364
rect 940 4336 948 4344
rect 1148 4336 1156 4344
rect 1388 4336 1396 4344
rect 1996 4336 2004 4344
rect 2076 4336 2084 4344
rect 2204 4336 2212 4344
rect 2268 4336 2276 4344
rect 2700 4336 2708 4344
rect 2908 4336 2916 4344
rect 3452 4336 3460 4344
rect 3532 4336 3540 4344
rect 4316 4336 4324 4344
rect 4460 4336 4468 4344
rect 4940 4336 4948 4344
rect 5708 4336 5716 4344
rect 5756 4336 5764 4344
rect 5964 4336 5972 4344
rect 6076 4336 6084 4344
rect 6124 4336 6132 4344
rect 6204 4336 6212 4344
rect 6748 4336 6756 4344
rect 6860 4336 6868 4344
rect 7196 4336 7204 4344
rect 7260 4336 7268 4344
rect 7420 4336 7428 4344
rect 7772 4336 7780 4344
rect 8092 4336 8100 4344
rect 60 4296 68 4304
rect 108 4316 116 4324
rect 300 4316 308 4324
rect 380 4316 388 4324
rect 428 4316 436 4324
rect 636 4316 644 4324
rect 700 4316 708 4324
rect 732 4316 740 4324
rect 972 4316 980 4324
rect 988 4316 996 4324
rect 1020 4316 1028 4324
rect 1052 4316 1060 4324
rect 1116 4316 1124 4324
rect 1260 4316 1268 4324
rect 1436 4316 1444 4324
rect 1500 4316 1508 4324
rect 1660 4316 1668 4324
rect 2028 4316 2036 4324
rect 2092 4316 2100 4324
rect 2156 4316 2164 4324
rect 2236 4316 2244 4324
rect 2396 4316 2404 4324
rect 2668 4316 2676 4324
rect 140 4296 148 4304
rect 172 4296 180 4304
rect 220 4296 228 4304
rect 284 4296 292 4304
rect 524 4296 532 4304
rect 92 4276 100 4284
rect 156 4276 164 4284
rect 28 4256 36 4264
rect 236 4276 244 4284
rect 332 4276 340 4284
rect 348 4276 356 4284
rect 476 4276 484 4284
rect 524 4276 532 4284
rect 636 4296 644 4304
rect 812 4296 820 4304
rect 1052 4296 1060 4304
rect 1100 4296 1108 4304
rect 1132 4296 1140 4304
rect 1180 4296 1188 4304
rect 1244 4296 1252 4304
rect 1292 4296 1300 4304
rect 1356 4296 1364 4304
rect 1404 4296 1412 4304
rect 1548 4296 1556 4304
rect 1628 4296 1636 4304
rect 1708 4296 1716 4304
rect 1772 4294 1780 4302
rect 1820 4296 1828 4304
rect 1916 4296 1924 4304
rect 1964 4296 1972 4304
rect 2012 4296 2020 4304
rect 2076 4296 2084 4304
rect 2204 4296 2212 4304
rect 2268 4296 2276 4304
rect 2364 4296 2372 4304
rect 2412 4296 2420 4304
rect 2460 4296 2468 4304
rect 2556 4296 2564 4304
rect 2700 4296 2708 4304
rect 2876 4316 2884 4324
rect 2940 4316 2948 4324
rect 3420 4316 3428 4324
rect 3836 4316 3844 4324
rect 2780 4296 2788 4304
rect 2812 4296 2820 4304
rect 2844 4296 2852 4304
rect 2924 4296 2932 4304
rect 2956 4296 2964 4304
rect 2988 4296 2996 4304
rect 3020 4296 3028 4304
rect 3132 4296 3140 4304
rect 3148 4296 3156 4304
rect 3292 4296 3300 4304
rect 3388 4296 3396 4304
rect 3436 4296 3444 4304
rect 3484 4296 3492 4304
rect 3660 4294 3668 4302
rect 3804 4296 3812 4304
rect 4012 4316 4020 4324
rect 4076 4316 4084 4324
rect 4284 4316 4292 4324
rect 4396 4316 4404 4324
rect 4428 4316 4436 4324
rect 4444 4316 4452 4324
rect 4588 4316 4596 4324
rect 4956 4316 4964 4324
rect 5148 4316 5156 4324
rect 3964 4296 3972 4304
rect 4076 4296 4084 4304
rect 4188 4296 4196 4304
rect 4316 4296 4324 4304
rect 4412 4296 4420 4304
rect 4476 4296 4484 4304
rect 4556 4296 4564 4304
rect 4588 4296 4596 4304
rect 4652 4294 4660 4302
rect 4716 4296 4724 4304
rect 4844 4296 4852 4304
rect 4892 4296 4900 4304
rect 4924 4296 4932 4304
rect 4988 4296 4996 4304
rect 5228 4296 5236 4304
rect 5260 4296 5268 4304
rect 5468 4296 5476 4304
rect 5500 4296 5508 4304
rect 5612 4296 5620 4304
rect 5708 4296 5716 4304
rect 6028 4316 6036 4324
rect 5788 4296 5796 4304
rect 5820 4296 5828 4304
rect 5884 4296 5892 4304
rect 5900 4296 5908 4304
rect 5996 4296 6004 4304
rect 6156 4316 6164 4324
rect 6172 4316 6180 4324
rect 6316 4316 6324 4324
rect 6348 4316 6356 4324
rect 6380 4316 6388 4324
rect 6460 4316 6468 4324
rect 6524 4316 6532 4324
rect 6828 4316 6836 4324
rect 7228 4316 7236 4324
rect 7244 4316 7252 4324
rect 7276 4316 7284 4324
rect 7324 4316 7332 4324
rect 7356 4316 7364 4324
rect 7388 4316 7396 4324
rect 7500 4316 7508 4324
rect 7596 4316 7604 4324
rect 7692 4316 7700 4324
rect 7740 4316 7748 4324
rect 6076 4296 6084 4304
rect 6140 4296 6148 4304
rect 6188 4296 6196 4304
rect 6236 4296 6244 4304
rect 6316 4296 6324 4304
rect 6700 4296 6708 4304
rect 684 4276 692 4284
rect 732 4276 740 4284
rect 780 4276 788 4284
rect 828 4276 836 4284
rect 940 4276 948 4284
rect 1036 4276 1044 4284
rect 1100 4276 1108 4284
rect 1196 4276 1204 4284
rect 1228 4276 1236 4284
rect 1244 4276 1252 4284
rect 1292 4276 1300 4284
rect 1404 4276 1412 4284
rect 1452 4276 1460 4284
rect 1532 4276 1540 4284
rect 1564 4280 1572 4288
rect 1612 4276 1620 4284
rect 1964 4276 1972 4284
rect 1996 4276 2004 4284
rect 2188 4276 2196 4284
rect 2252 4276 2260 4284
rect 2428 4276 2436 4284
rect 2572 4276 2580 4284
rect 2716 4276 2724 4284
rect 2764 4276 2772 4284
rect 2828 4276 2836 4284
rect 3628 4276 3636 4284
rect 3788 4276 3796 4284
rect 3804 4276 3812 4284
rect 3884 4276 3892 4284
rect 3916 4276 3924 4284
rect 3948 4276 3956 4284
rect 3980 4276 3988 4284
rect 4028 4276 4036 4284
rect 4172 4276 4180 4284
rect 4252 4276 4260 4284
rect 4620 4276 4628 4284
rect 4796 4276 4804 4284
rect 4972 4276 4980 4284
rect 5036 4276 5044 4284
rect 5132 4276 5140 4284
rect 5180 4276 5188 4284
rect 5244 4276 5252 4284
rect 5340 4276 5348 4284
rect 5356 4280 5364 4288
rect 5420 4276 5428 4284
rect 5596 4276 5604 4284
rect 5804 4276 5812 4284
rect 5836 4276 5844 4284
rect 5980 4276 5988 4284
rect 6092 4276 6100 4284
rect 6252 4276 6260 4284
rect 6300 4276 6308 4284
rect 6444 4276 6452 4284
rect 6492 4276 6500 4284
rect 6684 4276 6692 4284
rect 6716 4276 6724 4284
rect 6844 4296 6852 4304
rect 6908 4296 6916 4304
rect 7116 4294 7124 4302
rect 7212 4296 7220 4304
rect 7276 4296 7284 4304
rect 7324 4296 7332 4304
rect 7388 4296 7396 4304
rect 7500 4296 7508 4304
rect 7548 4296 7556 4304
rect 7580 4296 7588 4304
rect 7628 4296 7636 4304
rect 7788 4296 7796 4304
rect 7820 4296 7828 4304
rect 7900 4294 7908 4302
rect 8092 4296 8100 4304
rect 6892 4276 6900 4284
rect 6924 4276 6932 4284
rect 7148 4276 7156 4284
rect 7196 4276 7204 4284
rect 7308 4276 7316 4284
rect 7372 4276 7380 4284
rect 7452 4276 7460 4284
rect 7564 4276 7572 4284
rect 7772 4276 7780 4284
rect 7836 4276 7844 4284
rect 7916 4276 7924 4284
rect 8140 4276 8148 4284
rect 412 4256 420 4264
rect 444 4256 452 4264
rect 508 4256 516 4264
rect 636 4256 644 4264
rect 764 4256 772 4264
rect 1324 4256 1332 4264
rect 1516 4256 1524 4264
rect 1868 4256 1876 4264
rect 2108 4256 2116 4264
rect 2172 4256 2180 4264
rect 2316 4256 2324 4264
rect 2396 4256 2404 4264
rect 2460 4256 2468 4264
rect 2780 4256 2788 4264
rect 3020 4256 3028 4264
rect 3052 4256 3060 4264
rect 3260 4256 3268 4264
rect 3724 4256 3732 4264
rect 3756 4256 3764 4264
rect 4364 4256 4372 4264
rect 4508 4256 4516 4264
rect 5308 4256 5316 4264
rect 5660 4256 5668 4264
rect 5932 4256 5940 4264
rect 6204 4256 6212 4264
rect 6284 4256 6292 4264
rect 6412 4256 6420 4264
rect 6508 4256 6516 4264
rect 6572 4256 6580 4264
rect 6588 4256 6596 4264
rect 6620 4256 6628 4264
rect 6652 4256 6660 4264
rect 6956 4256 6964 4264
rect 7452 4256 7460 4264
rect 7676 4256 7684 4264
rect 7964 4256 7972 4264
rect 188 4236 196 4244
rect 252 4236 260 4244
rect 364 4236 372 4244
rect 492 4236 500 4244
rect 1196 4236 1204 4244
rect 1596 4236 1604 4244
rect 2476 4236 2484 4244
rect 2876 4236 2884 4244
rect 3068 4236 3076 4244
rect 4380 4236 4388 4244
rect 4780 4236 4788 4244
rect 5020 4236 5028 4244
rect 5068 4236 5076 4244
rect 5148 4236 5156 4244
rect 5196 4236 5204 4244
rect 5388 4236 5396 4244
rect 5644 4236 5652 4244
rect 5852 4236 5860 4244
rect 6268 4236 6276 4244
rect 6668 4236 6676 4244
rect 6844 4236 6852 4244
rect 6972 4236 6980 4244
rect 6988 4236 6996 4244
rect 7692 4236 7700 4244
rect 8044 4236 8052 4244
rect 8108 4236 8116 4244
rect 2172 4216 2180 4224
rect 2780 4216 2788 4224
rect 6508 4216 6516 4224
rect 3278 4206 3286 4214
rect 3292 4206 3300 4214
rect 3306 4206 3314 4214
rect 6350 4206 6358 4214
rect 6364 4206 6372 4214
rect 6378 4206 6386 4214
rect 556 4196 564 4204
rect 3052 4196 3060 4204
rect 6588 4196 6596 4204
rect 7548 4196 7556 4204
rect 76 4176 84 4184
rect 204 4176 212 4184
rect 508 4176 516 4184
rect 876 4176 884 4184
rect 1244 4176 1252 4184
rect 1532 4176 1540 4184
rect 1980 4176 1988 4184
rect 2012 4176 2020 4184
rect 2108 4176 2116 4184
rect 2540 4176 2548 4184
rect 2588 4176 2596 4184
rect 2668 4176 2676 4184
rect 2876 4176 2884 4184
rect 3020 4176 3028 4184
rect 3532 4176 3540 4184
rect 3756 4176 3764 4184
rect 3788 4176 3796 4184
rect 4044 4176 4052 4184
rect 4268 4176 4276 4184
rect 4700 4176 4708 4184
rect 4764 4176 4772 4184
rect 5244 4176 5252 4184
rect 5324 4176 5332 4184
rect 5468 4176 5476 4184
rect 5548 4176 5556 4184
rect 5596 4176 5604 4184
rect 5756 4176 5764 4184
rect 5788 4176 5796 4184
rect 6140 4176 6148 4184
rect 6188 4176 6196 4184
rect 6444 4176 6452 4184
rect 6972 4176 6980 4184
rect 7052 4176 7060 4184
rect 7116 4176 7124 4184
rect 7228 4176 7236 4184
rect 7292 4176 7300 4184
rect 7756 4176 7764 4184
rect 556 4156 564 4164
rect 620 4156 628 4164
rect 892 4156 900 4164
rect 908 4156 916 4164
rect 1020 4156 1028 4164
rect 1372 4156 1380 4164
rect 1724 4156 1732 4164
rect 1820 4156 1828 4164
rect 1996 4156 2004 4164
rect 12 4136 20 4144
rect 108 4136 116 4144
rect 140 4136 148 4144
rect 172 4136 180 4144
rect 236 4132 244 4140
rect 252 4136 260 4144
rect 476 4136 484 4144
rect 716 4136 724 4144
rect 860 4136 868 4144
rect 924 4136 932 4144
rect 1004 4136 1012 4144
rect 1084 4136 1092 4144
rect 1116 4136 1124 4144
rect 1436 4136 1444 4144
rect 1452 4132 1460 4140
rect 1500 4136 1508 4144
rect 1532 4136 1540 4144
rect 1580 4136 1588 4144
rect 1628 4136 1636 4144
rect 1868 4136 1876 4144
rect 1900 4136 1908 4144
rect 1932 4136 1940 4144
rect 2300 4156 2308 4164
rect 2492 4156 2500 4164
rect 2524 4156 2532 4164
rect 2684 4156 2692 4164
rect 2732 4156 2740 4164
rect 2044 4136 2052 4144
rect 2140 4136 2148 4144
rect 2188 4136 2196 4144
rect 28 4116 36 4124
rect 124 4116 132 4124
rect 188 4116 196 4124
rect 284 4116 292 4124
rect 428 4116 436 4124
rect 540 4116 548 4124
rect 652 4116 660 4124
rect 684 4116 692 4124
rect 748 4118 756 4126
rect 60 4096 68 4104
rect 76 4096 84 4104
rect 140 4096 148 4104
rect 268 4096 276 4104
rect 636 4096 644 4104
rect 956 4096 964 4104
rect 1036 4116 1044 4124
rect 1052 4116 1060 4124
rect 1068 4116 1076 4124
rect 1132 4116 1140 4124
rect 1164 4116 1172 4124
rect 1196 4116 1204 4124
rect 1356 4116 1364 4124
rect 1500 4116 1508 4124
rect 1644 4116 1652 4124
rect 1708 4116 1716 4124
rect 1756 4116 1764 4124
rect 1852 4116 1860 4124
rect 1916 4116 1924 4124
rect 2236 4116 2244 4124
rect 2332 4116 2340 4124
rect 2444 4116 2452 4124
rect 2508 4116 2516 4124
rect 2588 4116 2596 4124
rect 2812 4136 2820 4144
rect 2908 4136 2916 4144
rect 2988 4136 2996 4144
rect 3052 4156 3060 4164
rect 3116 4156 3124 4164
rect 3180 4156 3188 4164
rect 3356 4156 3364 4164
rect 3500 4156 3508 4164
rect 3772 4156 3780 4164
rect 4348 4156 4356 4164
rect 4412 4156 4420 4164
rect 4428 4156 4436 4164
rect 4492 4156 4500 4164
rect 4716 4156 4724 4164
rect 4780 4156 4788 4164
rect 4796 4156 4804 4164
rect 4860 4156 4868 4164
rect 5036 4156 5044 4164
rect 5116 4156 5124 4164
rect 5228 4156 5236 4164
rect 5308 4156 5316 4164
rect 5340 4156 5348 4164
rect 5660 4156 5668 4164
rect 5740 4156 5748 4164
rect 5772 4156 5780 4164
rect 6588 4156 6596 4164
rect 6652 4156 6660 4164
rect 7100 4156 7108 4164
rect 7164 4156 7172 4164
rect 7260 4156 7268 4164
rect 7308 4156 7316 4164
rect 7484 4156 7492 4164
rect 7548 4156 7556 4164
rect 7644 4156 7652 4164
rect 7708 4156 7716 4164
rect 8044 4156 8052 4164
rect 3052 4136 3060 4144
rect 3180 4136 3188 4144
rect 3212 4136 3220 4144
rect 3372 4136 3380 4144
rect 3468 4136 3476 4144
rect 3708 4136 3716 4144
rect 3804 4136 3812 4144
rect 3932 4136 3940 4144
rect 3996 4136 4004 4144
rect 4076 4136 4084 4144
rect 4108 4136 4116 4144
rect 4172 4136 4180 4144
rect 4316 4136 4324 4144
rect 4540 4136 4548 4144
rect 4700 4136 4708 4144
rect 4844 4136 4852 4144
rect 4972 4136 4980 4144
rect 5004 4136 5012 4144
rect 5148 4136 5156 4144
rect 5212 4136 5220 4144
rect 5292 4136 5300 4144
rect 2636 4116 2644 4124
rect 2716 4116 2724 4124
rect 2780 4116 2788 4124
rect 2956 4116 2964 4124
rect 2988 4116 2996 4124
rect 3132 4116 3140 4124
rect 3324 4116 3332 4124
rect 3468 4116 3476 4124
rect 3692 4116 3700 4124
rect 3724 4116 3732 4124
rect 3820 4116 3828 4124
rect 3900 4116 3908 4124
rect 3948 4116 3956 4124
rect 3964 4116 3972 4124
rect 1004 4096 1012 4104
rect 1116 4096 1124 4104
rect 1148 4096 1156 4104
rect 1532 4096 1540 4104
rect 1564 4096 1572 4104
rect 1628 4096 1636 4104
rect 1932 4096 1940 4104
rect 2156 4096 2164 4104
rect 2188 4096 2196 4104
rect 2604 4096 2612 4104
rect 2668 4096 2676 4104
rect 2700 4096 2708 4104
rect 2796 4096 2804 4104
rect 2972 4096 2980 4104
rect 3916 4096 3924 4104
rect 3980 4096 3988 4104
rect 4028 4096 4036 4104
rect 4156 4116 4164 4124
rect 4348 4116 4356 4124
rect 4492 4116 4500 4124
rect 4572 4116 4580 4124
rect 4716 4116 4724 4124
rect 4780 4116 4788 4124
rect 5052 4116 5060 4124
rect 5084 4116 5092 4124
rect 5116 4116 5124 4124
rect 5276 4116 5284 4124
rect 5372 4116 5380 4124
rect 5420 4116 5428 4124
rect 5452 4136 5460 4144
rect 5484 4136 5492 4144
rect 5516 4136 5524 4144
rect 5564 4136 5572 4144
rect 5644 4136 5652 4144
rect 5692 4136 5700 4144
rect 5740 4136 5748 4144
rect 5820 4136 5828 4144
rect 5852 4136 5860 4144
rect 6044 4136 6052 4144
rect 6076 4136 6084 4144
rect 6172 4136 6180 4144
rect 6252 4136 6260 4144
rect 6348 4136 6356 4144
rect 6460 4136 6468 4144
rect 6476 4136 6484 4144
rect 6524 4136 6532 4144
rect 6556 4136 6564 4144
rect 6732 4136 6740 4144
rect 6988 4136 6996 4144
rect 7084 4136 7092 4144
rect 7180 4136 7188 4144
rect 7196 4136 7204 4144
rect 7228 4136 7236 4144
rect 7276 4136 7284 4144
rect 7372 4136 7380 4144
rect 7388 4136 7396 4144
rect 7468 4136 7476 4144
rect 7708 4136 7716 4144
rect 7772 4136 7780 4144
rect 7788 4136 7796 4144
rect 7964 4136 7972 4144
rect 8012 4136 8020 4144
rect 8060 4136 8068 4144
rect 8092 4136 8100 4144
rect 5516 4116 5524 4124
rect 4316 4096 4324 4104
rect 4332 4096 4340 4104
rect 4508 4096 4516 4104
rect 4556 4096 4564 4104
rect 5100 4096 5108 4104
rect 5564 4096 5572 4104
rect 5836 4116 5844 4124
rect 5868 4116 5876 4124
rect 6012 4118 6020 4126
rect 6316 4118 6324 4126
rect 5612 4096 5620 4104
rect 5692 4096 5700 4104
rect 5724 4096 5732 4104
rect 6428 4096 6436 4104
rect 6508 4096 6516 4104
rect 6684 4116 6692 4124
rect 6748 4116 6756 4124
rect 6844 4118 6852 4126
rect 6892 4116 6900 4124
rect 7180 4116 7188 4124
rect 7244 4116 7252 4124
rect 7324 4116 7332 4124
rect 7356 4116 7364 4124
rect 6668 4096 6676 4104
rect 6748 4096 6756 4104
rect 6780 4096 6788 4104
rect 7308 4096 7316 4104
rect 7404 4096 7412 4104
rect 7548 4116 7556 4124
rect 7612 4116 7620 4124
rect 7660 4116 7668 4124
rect 7788 4116 7796 4124
rect 7884 4116 7892 4124
rect 7948 4116 7956 4124
rect 8140 4116 8148 4124
rect 7436 4096 7444 4104
rect 7836 4096 7844 4104
rect 7900 4096 7908 4104
rect 7980 4096 7988 4104
rect 668 4076 676 4084
rect 2572 4076 2580 4084
rect 2764 4076 2772 4084
rect 2940 4076 2948 4084
rect 3308 4076 3316 4084
rect 3884 4076 3892 4084
rect 4364 4076 4372 4084
rect 4540 4076 4548 4084
rect 2780 4056 2788 4064
rect 4588 4076 4596 4084
rect 4748 4076 4756 4084
rect 5036 4076 5044 4084
rect 5068 4076 5076 4084
rect 6620 4076 6628 4084
rect 6700 4076 6708 4084
rect 6940 4076 6948 4084
rect 7740 4076 7748 4084
rect 7868 4076 7876 4084
rect 6716 4056 6724 4064
rect 7900 4076 7908 4084
rect 8012 4076 8020 4084
rect 8092 4076 8100 4084
rect 28 4036 36 4044
rect 316 4036 324 4044
rect 588 4036 596 4044
rect 1692 4036 1700 4044
rect 1900 4036 1908 4044
rect 2428 4036 2436 4044
rect 2476 4036 2484 4044
rect 2540 4036 2548 4044
rect 2956 4036 2964 4044
rect 3084 4036 3092 4044
rect 3212 4036 3220 4044
rect 3420 4036 3428 4044
rect 3660 4036 3668 4044
rect 3820 4036 3828 4044
rect 4060 4036 4068 4044
rect 4396 4036 4404 4044
rect 4476 4036 4484 4044
rect 5324 4036 5332 4044
rect 5884 4036 5892 4044
rect 7356 4036 7364 4044
rect 7564 4036 7572 4044
rect 7804 4036 7812 4044
rect 7948 4036 7956 4044
rect 7996 4036 8004 4044
rect 1742 4006 1750 4014
rect 1756 4006 1764 4014
rect 1770 4006 1778 4014
rect 4814 4006 4822 4014
rect 4828 4006 4836 4014
rect 4842 4006 4850 4014
rect 12 3976 20 3984
rect 668 3976 676 3984
rect 732 3976 740 3984
rect 1164 3976 1172 3984
rect 1324 3976 1332 3984
rect 1372 3976 1380 3984
rect 1884 3976 1892 3984
rect 2380 3976 2388 3984
rect 2636 3976 2644 3984
rect 3052 3976 3060 3984
rect 3404 3976 3412 3984
rect 4348 3976 4356 3984
rect 4380 3976 4388 3984
rect 4412 3976 4420 3984
rect 4716 3976 4724 3984
rect 5228 3976 5236 3984
rect 5356 3976 5364 3984
rect 5612 3976 5620 3984
rect 7596 3976 7604 3984
rect 8044 3976 8052 3984
rect 8092 3976 8100 3984
rect 940 3956 948 3964
rect 3836 3956 3844 3964
rect 5852 3956 5860 3964
rect 7740 3956 7748 3964
rect 284 3936 292 3944
rect 476 3936 484 3944
rect 684 3936 692 3944
rect 1388 3936 1396 3944
rect 2316 3936 2324 3944
rect 3868 3936 3876 3944
rect 4364 3936 4372 3944
rect 4684 3936 4692 3944
rect 4732 3936 4740 3944
rect 4892 3936 4900 3944
rect 4956 3936 4964 3944
rect 5340 3936 5348 3944
rect 5372 3936 5380 3944
rect 5868 3936 5876 3944
rect 5948 3936 5956 3944
rect 6668 3936 6676 3944
rect 6860 3936 6868 3944
rect 8108 3936 8116 3944
rect 588 3916 596 3924
rect 652 3916 660 3924
rect 92 3894 100 3902
rect 412 3894 420 3902
rect 524 3896 532 3904
rect 556 3896 564 3904
rect 620 3896 628 3904
rect 668 3896 676 3904
rect 732 3896 740 3904
rect 780 3916 788 3924
rect 844 3916 852 3924
rect 1052 3916 1060 3924
rect 812 3896 820 3904
rect 876 3896 884 3904
rect 1628 3916 1636 3924
rect 1868 3916 1876 3924
rect 1932 3916 1940 3924
rect 2300 3916 2308 3924
rect 2412 3916 2420 3924
rect 2508 3916 2516 3924
rect 2700 3916 2708 3924
rect 2732 3916 2740 3924
rect 3084 3916 3092 3924
rect 3372 3916 3380 3924
rect 3548 3916 3556 3924
rect 3628 3916 3636 3924
rect 3708 3916 3716 3924
rect 3740 3916 3748 3924
rect 3772 3916 3780 3924
rect 4060 3916 4068 3924
rect 4396 3916 4404 3924
rect 4652 3916 4660 3924
rect 5196 3916 5204 3924
rect 5324 3916 5332 3924
rect 5708 3916 5716 3924
rect 5740 3916 5748 3924
rect 5804 3916 5812 3924
rect 5820 3916 5828 3924
rect 5900 3916 5908 3924
rect 6204 3916 6212 3924
rect 6620 3916 6628 3924
rect 6876 3916 6884 3924
rect 6908 3916 6916 3924
rect 7356 3916 7364 3924
rect 7372 3916 7380 3924
rect 7612 3916 7620 3924
rect 8012 3916 8020 3924
rect 8076 3916 8084 3924
rect 1148 3896 1156 3904
rect 1276 3896 1284 3904
rect 1420 3896 1428 3904
rect 1516 3896 1524 3904
rect 1628 3896 1636 3904
rect 1660 3896 1668 3904
rect 1804 3896 1812 3904
rect 1868 3896 1876 3904
rect 1964 3896 1972 3904
rect 2092 3896 2100 3904
rect 2268 3896 2276 3904
rect 2284 3896 2292 3904
rect 2380 3896 2388 3904
rect 2428 3896 2436 3904
rect 2508 3896 2516 3904
rect 2524 3896 2532 3904
rect 2540 3896 2548 3904
rect 2572 3896 2580 3904
rect 2604 3896 2612 3904
rect 2684 3896 2692 3904
rect 2956 3896 2964 3904
rect 3052 3896 3060 3904
rect 3148 3894 3156 3902
rect 3196 3896 3204 3904
rect 3388 3896 3396 3904
rect 3452 3896 3460 3904
rect 3468 3896 3476 3904
rect 3500 3896 3508 3904
rect 3580 3896 3588 3904
rect 3660 3896 3668 3904
rect 3724 3896 3732 3904
rect 3740 3896 3748 3904
rect 3788 3896 3796 3904
rect 3852 3896 3860 3904
rect 3932 3896 3940 3904
rect 3980 3896 3988 3904
rect 4076 3896 4084 3904
rect 4092 3896 4100 3904
rect 4204 3894 4212 3902
rect 4380 3896 4388 3904
rect 4444 3896 4452 3904
rect 4508 3894 4516 3902
rect 4668 3896 4676 3904
rect 4748 3896 4756 3904
rect 4940 3896 4948 3904
rect 5196 3896 5204 3904
rect 5228 3896 5236 3904
rect 5260 3896 5268 3904
rect 5324 3896 5332 3904
rect 5532 3896 5540 3904
rect 5644 3896 5652 3904
rect 5740 3896 5748 3904
rect 5788 3896 5796 3904
rect 5852 3896 5860 3904
rect 6060 3894 6068 3902
rect 6220 3896 6228 3904
rect 6236 3896 6244 3904
rect 6396 3894 6404 3902
rect 6588 3896 6596 3904
rect 6716 3896 6724 3904
rect 6828 3896 6836 3904
rect 6908 3896 6916 3904
rect 7084 3896 7092 3904
rect 7324 3896 7332 3904
rect 7356 3896 7364 3904
rect 7468 3894 7476 3902
rect 7692 3896 7700 3904
rect 7868 3896 7876 3904
rect 7948 3896 7956 3904
rect 7996 3896 8004 3904
rect 8044 3896 8052 3904
rect 124 3876 132 3884
rect 236 3876 244 3884
rect 508 3876 516 3884
rect 540 3876 548 3884
rect 636 3876 644 3884
rect 716 3876 724 3884
rect 828 3876 836 3884
rect 908 3876 916 3884
rect 1004 3876 1012 3884
rect 1020 3876 1028 3884
rect 1100 3876 1108 3884
rect 1196 3880 1204 3888
rect 1212 3876 1220 3884
rect 1260 3876 1268 3884
rect 1452 3876 1460 3884
rect 1820 3876 1828 3884
rect 2044 3876 2052 3884
rect 2348 3876 2356 3884
rect 2364 3876 2372 3884
rect 2444 3876 2452 3884
rect 2460 3876 2468 3884
rect 2492 3876 2500 3884
rect 2556 3876 2564 3884
rect 2636 3876 2644 3884
rect 2668 3876 2676 3884
rect 2684 3876 2692 3884
rect 2732 3876 2740 3884
rect 2796 3876 2804 3884
rect 2828 3876 2836 3884
rect 3004 3876 3012 3884
rect 3036 3876 3044 3884
rect 3116 3876 3124 3884
rect 3340 3876 3348 3884
rect 3436 3876 3444 3884
rect 28 3856 36 3864
rect 412 3856 420 3864
rect 860 3856 868 3864
rect 892 3856 900 3864
rect 1244 3856 1252 3864
rect 1356 3856 1364 3864
rect 1756 3856 1764 3864
rect 1852 3856 1860 3864
rect 1916 3856 1924 3864
rect 2012 3856 2020 3864
rect 2572 3856 2580 3864
rect 2604 3856 2612 3864
rect 2748 3856 2756 3864
rect 2828 3856 2836 3864
rect 3516 3876 3524 3884
rect 3564 3876 3572 3884
rect 3724 3876 3732 3884
rect 3804 3876 3812 3884
rect 3836 3876 3844 3884
rect 4028 3876 4036 3884
rect 4172 3876 4180 3884
rect 4476 3876 4484 3884
rect 4860 3876 4868 3884
rect 4988 3876 4996 3884
rect 5132 3876 5140 3884
rect 5148 3880 5156 3888
rect 5404 3876 5412 3884
rect 5452 3876 5460 3884
rect 5500 3876 5508 3884
rect 5628 3876 5636 3884
rect 5692 3876 5700 3884
rect 5932 3876 5940 3884
rect 5980 3876 5988 3884
rect 6364 3876 6372 3884
rect 6620 3876 6628 3884
rect 6796 3876 6804 3884
rect 7132 3876 7140 3884
rect 7164 3876 7172 3884
rect 7292 3876 7300 3884
rect 7308 3876 7316 3884
rect 7372 3876 7380 3884
rect 7404 3876 7412 3884
rect 7484 3876 7492 3884
rect 7644 3876 7652 3884
rect 7708 3876 7716 3884
rect 7916 3876 7924 3884
rect 7980 3876 7988 3884
rect 8092 3896 8100 3904
rect 3628 3856 3636 3864
rect 4140 3856 4148 3864
rect 4796 3856 4804 3864
rect 4876 3856 4884 3864
rect 4972 3856 4980 3864
rect 5292 3856 5300 3864
rect 5420 3856 5428 3864
rect 5756 3856 5764 3864
rect 5820 3856 5828 3864
rect 5900 3856 5908 3864
rect 5996 3856 6004 3864
rect 6060 3856 6068 3864
rect 6284 3856 6292 3864
rect 6540 3856 6548 3864
rect 7724 3856 7732 3864
rect 7948 3856 7956 3864
rect 220 3836 228 3844
rect 252 3836 260 3844
rect 492 3836 500 3844
rect 1068 3836 1076 3844
rect 1116 3836 1124 3844
rect 1612 3836 1620 3844
rect 1724 3836 1732 3844
rect 1932 3836 1940 3844
rect 2204 3836 2212 3844
rect 2316 3836 2324 3844
rect 2844 3836 2852 3844
rect 3276 3836 3284 3844
rect 3548 3836 3556 3844
rect 4332 3836 4340 3844
rect 4636 3836 4644 3844
rect 4668 3836 4676 3844
rect 4924 3836 4932 3844
rect 5100 3836 5108 3844
rect 6188 3836 6196 3844
rect 6524 3836 6532 3844
rect 6636 3836 6644 3844
rect 6972 3836 6980 3844
rect 7612 3836 7620 3844
rect 7660 3836 7668 3844
rect 7756 3836 7764 3844
rect 3278 3806 3286 3814
rect 3292 3806 3300 3814
rect 3306 3806 3314 3814
rect 6350 3806 6358 3814
rect 6364 3806 6372 3814
rect 6378 3806 6386 3814
rect 4284 3796 4292 3804
rect 6172 3796 6180 3804
rect 188 3776 196 3784
rect 620 3776 628 3784
rect 700 3776 708 3784
rect 1436 3776 1444 3784
rect 1580 3776 1588 3784
rect 1852 3776 1860 3784
rect 1884 3776 1892 3784
rect 2092 3776 2100 3784
rect 2252 3776 2260 3784
rect 2364 3776 2372 3784
rect 2396 3776 2404 3784
rect 2492 3776 2500 3784
rect 2524 3776 2532 3784
rect 2732 3776 2740 3784
rect 2940 3776 2948 3784
rect 2972 3776 2980 3784
rect 3180 3776 3188 3784
rect 3212 3776 3220 3784
rect 3644 3776 3652 3784
rect 3724 3776 3732 3784
rect 4204 3776 4212 3784
rect 4428 3776 4436 3784
rect 4972 3776 4980 3784
rect 5388 3776 5396 3784
rect 5532 3776 5540 3784
rect 5788 3776 5796 3784
rect 5868 3776 5876 3784
rect 6028 3776 6036 3784
rect 6492 3776 6500 3784
rect 6556 3776 6564 3784
rect 6668 3776 6676 3784
rect 6684 3776 6692 3784
rect 6860 3776 6868 3784
rect 6908 3776 6916 3784
rect 7180 3776 7188 3784
rect 8108 3776 8116 3784
rect 204 3756 212 3764
rect 572 3756 580 3764
rect 588 3756 596 3764
rect 892 3756 900 3764
rect 924 3756 932 3764
rect 1068 3756 1076 3764
rect 1244 3756 1252 3764
rect 1308 3756 1316 3764
rect 1468 3756 1476 3764
rect 1516 3756 1524 3764
rect 1740 3756 1748 3764
rect 1900 3756 1908 3764
rect 1964 3756 1972 3764
rect 2140 3756 2148 3764
rect 2268 3756 2276 3764
rect 2316 3756 2324 3764
rect 2380 3756 2388 3764
rect 2924 3756 2932 3764
rect 3052 3756 3060 3764
rect 3196 3756 3204 3764
rect 3484 3756 3492 3764
rect 3500 3756 3508 3764
rect 3676 3756 3684 3764
rect 3708 3756 3716 3764
rect 3788 3756 3796 3764
rect 4012 3756 4020 3764
rect 4220 3756 4228 3764
rect 4284 3756 4292 3764
rect 4300 3756 4308 3764
rect 4396 3756 4404 3764
rect 4556 3756 4564 3764
rect 4716 3756 4724 3764
rect 4748 3756 4756 3764
rect 4828 3756 4836 3764
rect 4956 3756 4964 3764
rect 5052 3756 5060 3764
rect 5260 3756 5268 3764
rect 5420 3756 5428 3764
rect 5452 3756 5460 3764
rect 5836 3756 5844 3764
rect 6124 3756 6132 3764
rect 6172 3756 6180 3764
rect 6236 3756 6244 3764
rect 6588 3756 6596 3764
rect 316 3736 324 3744
rect 492 3736 500 3744
rect 540 3736 548 3744
rect 572 3736 580 3744
rect 652 3736 660 3744
rect 668 3736 676 3744
rect 700 3736 708 3744
rect 732 3736 740 3744
rect 764 3736 772 3744
rect 796 3736 804 3744
rect 956 3736 964 3744
rect 1020 3732 1028 3740
rect 1036 3736 1044 3744
rect 1084 3736 1092 3744
rect 1100 3736 1108 3744
rect 1196 3736 1204 3744
rect 1484 3736 1492 3744
rect 1532 3736 1540 3744
rect 1612 3736 1620 3744
rect 1644 3736 1652 3744
rect 1708 3736 1716 3744
rect 1804 3736 1812 3744
rect 2108 3736 2116 3744
rect 2156 3736 2164 3744
rect 2220 3736 2228 3744
rect 2284 3736 2292 3744
rect 2348 3736 2356 3744
rect 2444 3736 2452 3744
rect 2508 3736 2516 3744
rect 2588 3736 2596 3744
rect 2652 3736 2660 3744
rect 2684 3736 2692 3744
rect 2780 3736 2788 3744
rect 2796 3736 2804 3744
rect 2844 3736 2852 3744
rect 2876 3736 2884 3744
rect 2908 3736 2916 3744
rect 2988 3736 2996 3744
rect 3276 3736 3284 3744
rect 3452 3736 3460 3744
rect 3468 3736 3476 3744
rect 3516 3736 3524 3744
rect 3532 3736 3540 3744
rect 3564 3736 3572 3744
rect 3596 3736 3604 3744
rect 3708 3736 3716 3744
rect 3948 3736 3956 3744
rect 4108 3736 4116 3744
rect 4412 3736 4420 3744
rect 4620 3736 4628 3744
rect 4652 3736 4660 3744
rect 4732 3736 4740 3744
rect 4812 3736 4820 3744
rect 5068 3736 5076 3744
rect 5436 3736 5444 3744
rect 5708 3736 5716 3744
rect 5788 3736 5796 3744
rect 5836 3736 5844 3744
rect 5852 3736 5860 3744
rect 5916 3736 5924 3744
rect 5980 3736 5988 3744
rect 6060 3736 6068 3744
rect 6156 3736 6164 3744
rect 6252 3736 6260 3744
rect 6268 3732 6276 3740
rect 6316 3736 6324 3744
rect 6428 3736 6436 3744
rect 6444 3736 6452 3744
rect 6460 3736 6468 3744
rect 6492 3736 6500 3744
rect 6748 3736 6756 3744
rect 7372 3756 7380 3764
rect 7596 3756 7604 3764
rect 7692 3756 7700 3764
rect 6780 3736 6788 3744
rect 6876 3736 6884 3744
rect 6940 3736 6948 3744
rect 7148 3736 7156 3744
rect 7340 3736 7348 3744
rect 7436 3736 7444 3744
rect 7468 3736 7476 3744
rect 7532 3736 7540 3744
rect 7548 3736 7556 3744
rect 7676 3736 7684 3744
rect 7772 3736 7780 3744
rect 7868 3736 7876 3744
rect 7900 3736 7908 3744
rect 7916 3736 7924 3744
rect 7948 3736 7956 3744
rect 92 3716 100 3724
rect 124 3716 132 3724
rect 252 3716 260 3724
rect 268 3716 276 3724
rect 348 3718 356 3726
rect 412 3716 420 3724
rect 524 3716 532 3724
rect 716 3716 724 3724
rect 780 3716 788 3724
rect 812 3716 820 3724
rect 844 3716 852 3724
rect 908 3716 916 3724
rect 972 3716 980 3724
rect 988 3716 996 3724
rect 1116 3716 1124 3724
rect 1212 3716 1220 3724
rect 1308 3718 1316 3726
rect 1484 3716 1492 3724
rect 1532 3716 1540 3724
rect 1548 3716 1556 3724
rect 156 3696 164 3704
rect 284 3696 292 3704
rect 700 3696 708 3704
rect 844 3696 852 3704
rect 1596 3716 1604 3724
rect 1820 3716 1828 3724
rect 1868 3716 1876 3724
rect 1964 3718 1972 3726
rect 2140 3716 2148 3724
rect 2220 3716 2228 3724
rect 2300 3716 2308 3724
rect 2460 3716 2468 3724
rect 1676 3696 1684 3704
rect 2204 3696 2212 3704
rect 2252 3696 2260 3704
rect 2396 3696 2404 3704
rect 2604 3716 2612 3724
rect 2684 3716 2692 3724
rect 2812 3716 2820 3724
rect 2556 3696 2564 3704
rect 2860 3716 2868 3724
rect 2892 3716 2900 3724
rect 3052 3718 3060 3726
rect 3276 3716 3284 3724
rect 3356 3716 3364 3724
rect 3436 3716 3444 3724
rect 3548 3716 3556 3724
rect 3788 3718 3796 3726
rect 3980 3716 3988 3724
rect 4076 3718 4084 3726
rect 4364 3716 4372 3724
rect 4396 3716 4404 3724
rect 4556 3718 4564 3726
rect 4620 3716 4628 3724
rect 4668 3716 4676 3724
rect 4828 3716 4836 3724
rect 4908 3716 4916 3724
rect 4924 3716 4932 3724
rect 2860 3696 2868 3704
rect 2956 3696 2964 3704
rect 3228 3696 3236 3704
rect 3340 3696 3348 3704
rect 3404 3696 3412 3704
rect 3644 3696 3652 3704
rect 3660 3696 3668 3704
rect 3932 3696 3940 3704
rect 4668 3696 4676 3704
rect 4764 3696 4772 3704
rect 4780 3696 4788 3704
rect 4892 3696 4900 3704
rect 5020 3716 5028 3724
rect 5196 3716 5204 3724
rect 5260 3718 5268 3726
rect 5500 3716 5508 3724
rect 5612 3716 5620 3724
rect 5676 3718 5684 3726
rect 5740 3716 5748 3724
rect 5900 3716 5908 3724
rect 5964 3716 5972 3724
rect 6076 3716 6084 3724
rect 6156 3716 6164 3724
rect 6300 3716 6308 3724
rect 5404 3696 5412 3704
rect 5532 3696 5540 3704
rect 5788 3696 5796 3704
rect 5932 3696 5940 3704
rect 6028 3696 6036 3704
rect 6044 3696 6052 3704
rect 6108 3696 6116 3704
rect 6124 3696 6132 3704
rect 6396 3696 6404 3704
rect 6508 3716 6516 3724
rect 6572 3716 6580 3724
rect 6620 3716 6628 3724
rect 6636 3716 6644 3724
rect 6732 3716 6740 3724
rect 6828 3716 6836 3724
rect 6892 3716 6900 3724
rect 7116 3718 7124 3726
rect 7308 3718 7316 3726
rect 7420 3716 7428 3724
rect 7580 3716 7588 3724
rect 7628 3716 7636 3724
rect 7692 3716 7700 3724
rect 7724 3716 7732 3724
rect 6492 3696 6500 3704
rect 6812 3696 6820 3704
rect 7452 3696 7460 3704
rect 7500 3696 7508 3704
rect 7644 3696 7652 3704
rect 7820 3716 7828 3724
rect 7836 3716 7844 3724
rect 7916 3716 7924 3724
rect 7980 3718 7988 3726
rect 8044 3716 8052 3724
rect 492 3676 500 3684
rect 1036 3676 1044 3684
rect 2316 3676 2324 3684
rect 3196 3676 3204 3684
rect 3372 3676 3380 3684
rect 3612 3676 3620 3684
rect 3916 3676 3924 3684
rect 6044 3676 6052 3684
rect 6684 3676 6692 3684
rect 6908 3676 6916 3684
rect 6988 3676 6996 3684
rect 7788 3676 7796 3684
rect 7900 3676 7908 3684
rect 764 3656 772 3664
rect 1724 3656 1732 3664
rect 3260 3656 3268 3664
rect 812 3636 820 3644
rect 1436 3636 1444 3644
rect 1452 3636 1460 3644
rect 1612 3636 1620 3644
rect 2668 3636 2676 3644
rect 3356 3636 3364 3644
rect 3436 3636 3444 3644
rect 3580 3636 3588 3644
rect 4252 3636 4260 3644
rect 4316 3636 4324 3644
rect 4332 3636 4340 3644
rect 4684 3636 4692 3644
rect 5548 3636 5556 3644
rect 5964 3636 5972 3644
rect 6076 3636 6084 3644
rect 6956 3636 6964 3644
rect 1742 3606 1750 3614
rect 1756 3606 1764 3614
rect 1770 3606 1778 3614
rect 4814 3606 4822 3614
rect 4828 3606 4836 3614
rect 4842 3606 4850 3614
rect 92 3576 100 3584
rect 940 3576 948 3584
rect 1308 3576 1316 3584
rect 1580 3576 1588 3584
rect 2012 3576 2020 3584
rect 2028 3576 2036 3584
rect 2988 3576 2996 3584
rect 3036 3576 3044 3584
rect 3452 3576 3460 3584
rect 4508 3576 4516 3584
rect 4636 3576 4644 3584
rect 4940 3576 4948 3584
rect 5260 3576 5268 3584
rect 5436 3576 5444 3584
rect 5788 3576 5796 3584
rect 6284 3576 6292 3584
rect 6828 3576 6836 3584
rect 7164 3576 7172 3584
rect 7308 3576 7316 3584
rect 7788 3576 7796 3584
rect 8092 3576 8100 3584
rect 1100 3556 1108 3564
rect 3804 3556 3812 3564
rect 5340 3556 5348 3564
rect 7004 3556 7012 3564
rect 108 3536 116 3544
rect 1292 3536 1300 3544
rect 1372 3536 1380 3544
rect 1404 3536 1412 3544
rect 2652 3536 2660 3544
rect 2972 3536 2980 3544
rect 3244 3536 3252 3544
rect 3628 3536 3636 3544
rect 3852 3536 3860 3544
rect 4268 3536 4276 3544
rect 4524 3536 4532 3544
rect 5084 3536 5092 3544
rect 5324 3536 5332 3544
rect 5724 3536 5732 3544
rect 5804 3536 5812 3544
rect 5900 3536 5908 3544
rect 6300 3536 6308 3544
rect 6380 3536 6388 3544
rect 6524 3536 6532 3544
rect 6620 3536 6628 3544
rect 6860 3536 6868 3544
rect 7180 3536 7188 3544
rect 7244 3536 7252 3544
rect 7324 3536 7332 3544
rect 12 3516 20 3524
rect 76 3516 84 3524
rect 188 3516 196 3524
rect 268 3516 276 3524
rect 492 3516 500 3524
rect 1052 3516 1060 3524
rect 44 3496 52 3504
rect 92 3496 100 3504
rect 332 3496 340 3504
rect 460 3496 468 3504
rect 524 3496 532 3504
rect 620 3496 628 3504
rect 668 3496 676 3504
rect 812 3496 820 3504
rect 860 3496 868 3504
rect 1004 3496 1012 3504
rect 1132 3516 1140 3524
rect 1228 3516 1236 3524
rect 1324 3516 1332 3524
rect 1340 3516 1348 3524
rect 1516 3516 1524 3524
rect 1596 3516 1604 3524
rect 2268 3516 2276 3524
rect 2300 3516 2308 3524
rect 2348 3516 2356 3524
rect 1228 3496 1236 3504
rect 1308 3496 1316 3504
rect 1356 3496 1364 3504
rect 1436 3496 1444 3504
rect 1500 3496 1508 3504
rect 1628 3496 1636 3504
rect 1660 3496 1668 3504
rect 1676 3496 1684 3504
rect 1884 3494 1892 3502
rect 2156 3494 2164 3502
rect 2268 3496 2276 3504
rect 2556 3516 2564 3524
rect 2620 3516 2628 3524
rect 2748 3516 2756 3524
rect 2796 3516 2804 3524
rect 2860 3516 2868 3524
rect 2940 3516 2948 3524
rect 3004 3516 3012 3524
rect 3052 3516 3060 3524
rect 3356 3516 3364 3524
rect 3388 3516 3396 3524
rect 3420 3516 3428 3524
rect 3596 3516 3604 3524
rect 3660 3516 3668 3524
rect 3772 3516 3780 3524
rect 3884 3516 3892 3524
rect 4380 3516 4388 3524
rect 4444 3516 4452 3524
rect 4492 3516 4500 3524
rect 4556 3516 4564 3524
rect 2476 3496 2484 3504
rect 2540 3496 2548 3504
rect 2604 3496 2612 3504
rect 2716 3496 2724 3504
rect 2908 3496 2916 3504
rect 2924 3496 2932 3504
rect 2988 3496 2996 3504
rect 3132 3496 3140 3504
rect 3436 3496 3444 3504
rect 3500 3496 3508 3504
rect 3644 3496 3652 3504
rect 3692 3496 3700 3504
rect 3740 3496 3748 3504
rect 3772 3496 3780 3504
rect 3804 3496 3812 3504
rect 3868 3496 3876 3504
rect 3996 3496 4004 3504
rect 4156 3496 4164 3504
rect 4284 3496 4292 3504
rect 4332 3496 4340 3504
rect 4364 3496 4372 3504
rect 4508 3496 4516 3504
rect 4556 3496 4564 3504
rect 4604 3496 4612 3504
rect 4620 3496 4628 3504
rect 4748 3516 4756 3524
rect 4972 3516 4980 3524
rect 5004 3516 5012 3524
rect 5356 3516 5364 3524
rect 5372 3516 5380 3524
rect 5612 3516 5620 3524
rect 5644 3516 5652 3524
rect 5660 3516 5668 3524
rect 5756 3516 5764 3524
rect 5772 3516 5780 3524
rect 5852 3516 5860 3524
rect 6268 3516 6276 3524
rect 6332 3516 6340 3524
rect 6604 3516 6612 3524
rect 6892 3516 6900 3524
rect 6956 3516 6964 3524
rect 4828 3496 4836 3504
rect 4892 3496 4900 3504
rect 4956 3496 4964 3504
rect 5196 3496 5204 3504
rect 5212 3496 5220 3504
rect 5292 3496 5300 3504
rect 5340 3496 5348 3504
rect 5420 3496 5428 3504
rect 5484 3496 5492 3504
rect 5500 3496 5508 3504
rect 5548 3496 5556 3504
rect 5612 3496 5620 3504
rect 5644 3496 5652 3504
rect 5692 3496 5700 3504
rect 5788 3496 5796 3504
rect 5948 3496 5956 3504
rect 6012 3496 6020 3504
rect 6092 3496 6100 3504
rect 6108 3496 6116 3504
rect 6172 3496 6180 3504
rect 6188 3496 6196 3504
rect 6252 3496 6260 3504
rect 6284 3496 6292 3504
rect 6476 3496 6484 3504
rect 6572 3496 6580 3504
rect 6716 3496 6724 3504
rect 6876 3496 6884 3504
rect 6924 3496 6932 3504
rect 7020 3496 7028 3504
rect 7148 3516 7156 3524
rect 7724 3516 7732 3524
rect 7164 3496 7172 3504
rect 7436 3496 7444 3504
rect 7516 3496 7524 3504
rect 7900 3496 7908 3504
rect 60 3476 68 3484
rect 140 3476 148 3484
rect 156 3456 164 3464
rect 172 3456 180 3464
rect 236 3456 244 3464
rect 252 3456 260 3464
rect 316 3456 324 3464
rect 364 3456 372 3464
rect 476 3476 484 3484
rect 540 3476 548 3484
rect 572 3476 580 3484
rect 1004 3476 1012 3484
rect 1116 3476 1124 3484
rect 1164 3476 1172 3484
rect 1180 3476 1188 3484
rect 1372 3476 1380 3484
rect 1452 3476 1460 3484
rect 1548 3476 1556 3484
rect 1564 3476 1572 3484
rect 1644 3476 1652 3484
rect 1676 3476 1684 3484
rect 1788 3476 1796 3484
rect 2140 3476 2148 3484
rect 2316 3476 2324 3484
rect 2396 3476 2404 3484
rect 2428 3476 2436 3484
rect 2444 3476 2452 3484
rect 2556 3476 2564 3484
rect 2588 3476 2596 3484
rect 2604 3476 2612 3484
rect 956 3456 964 3464
rect 972 3456 980 3464
rect 1260 3456 1268 3464
rect 1420 3456 1428 3464
rect 1612 3456 1620 3464
rect 1884 3456 1892 3464
rect 2764 3476 2772 3484
rect 2892 3476 2900 3484
rect 3020 3476 3028 3484
rect 3260 3476 3268 3484
rect 3388 3476 3396 3484
rect 3484 3476 3492 3484
rect 3516 3476 3524 3484
rect 3564 3476 3572 3484
rect 3628 3476 3636 3484
rect 3676 3476 3684 3484
rect 3820 3476 3828 3484
rect 3868 3476 3876 3484
rect 4060 3476 4068 3484
rect 4108 3476 4116 3484
rect 4364 3476 4372 3484
rect 4428 3476 4436 3484
rect 4476 3476 4484 3484
rect 4620 3476 4628 3484
rect 4636 3476 4644 3484
rect 4668 3476 4676 3484
rect 4700 3476 4708 3484
rect 4796 3476 4804 3484
rect 4812 3476 4820 3484
rect 4908 3476 4916 3484
rect 5004 3476 5012 3484
rect 5036 3476 5044 3484
rect 5100 3476 5108 3484
rect 5196 3476 5204 3484
rect 5228 3476 5236 3484
rect 5404 3476 5412 3484
rect 5436 3476 5444 3484
rect 5468 3476 5476 3484
rect 5500 3476 5508 3484
rect 5692 3476 5700 3484
rect 5980 3476 5988 3484
rect 5996 3476 6004 3484
rect 6124 3476 6132 3484
rect 6156 3476 6164 3484
rect 6204 3476 6212 3484
rect 6236 3476 6244 3484
rect 6364 3476 6372 3484
rect 6508 3476 6516 3484
rect 6604 3476 6612 3484
rect 6876 3476 6884 3484
rect 6908 3476 6916 3484
rect 7020 3476 7028 3484
rect 7068 3476 7076 3484
rect 7084 3476 7092 3484
rect 7484 3476 7492 3484
rect 7644 3476 7652 3484
rect 7692 3476 7700 3484
rect 7772 3476 7780 3484
rect 7948 3476 7956 3484
rect 7980 3476 7988 3484
rect 2092 3456 2100 3464
rect 2220 3456 2228 3464
rect 2492 3456 2500 3464
rect 2668 3456 2676 3464
rect 2812 3456 2820 3464
rect 2876 3456 2884 3464
rect 3116 3456 3124 3464
rect 3356 3456 3364 3464
rect 3740 3456 3748 3464
rect 4332 3456 4340 3464
rect 4364 3456 4372 3464
rect 4796 3456 4804 3464
rect 5036 3456 5044 3464
rect 5260 3456 5268 3464
rect 5276 3456 5284 3464
rect 5580 3456 5588 3464
rect 5836 3456 5844 3464
rect 5900 3456 5908 3464
rect 5932 3456 5940 3464
rect 6060 3456 6068 3464
rect 6092 3456 6100 3464
rect 6332 3456 6340 3464
rect 6444 3456 6452 3464
rect 6524 3456 6532 3464
rect 6748 3456 6756 3464
rect 6812 3456 6820 3464
rect 7212 3456 7220 3464
rect 7276 3456 7284 3464
rect 7292 3456 7300 3464
rect 7660 3456 7668 3464
rect 12 3436 20 3444
rect 396 3436 404 3444
rect 492 3436 500 3444
rect 732 3436 740 3444
rect 924 3436 932 3444
rect 988 3436 996 3444
rect 1228 3436 1236 3444
rect 1484 3436 1492 3444
rect 2012 3436 2020 3444
rect 2748 3436 2756 3444
rect 2796 3436 2804 3444
rect 3340 3436 3348 3444
rect 3532 3436 3540 3444
rect 3900 3436 3908 3444
rect 5020 3436 5028 3444
rect 5068 3436 5076 3444
rect 5388 3436 5396 3444
rect 6044 3436 6052 3444
rect 6156 3436 6164 3444
rect 6220 3436 6228 3444
rect 7132 3436 7140 3444
rect 7676 3436 7684 3444
rect 7756 3436 7764 3444
rect 172 3416 180 3424
rect 252 3416 260 3424
rect 2876 3416 2884 3424
rect 4364 3416 4372 3424
rect 5836 3416 5844 3424
rect 3278 3406 3286 3414
rect 3292 3406 3300 3414
rect 3306 3406 3314 3414
rect 6350 3406 6358 3414
rect 6364 3406 6372 3414
rect 6378 3406 6386 3414
rect 1388 3396 1396 3404
rect 1756 3396 1764 3404
rect 2828 3396 2836 3404
rect 7148 3396 7156 3404
rect 7276 3396 7284 3404
rect 92 3376 100 3384
rect 140 3376 148 3384
rect 236 3376 244 3384
rect 492 3376 500 3384
rect 1260 3376 1268 3384
rect 1740 3376 1748 3384
rect 1948 3376 1956 3384
rect 2172 3376 2180 3384
rect 2940 3376 2948 3384
rect 3004 3376 3012 3384
rect 3340 3376 3348 3384
rect 3500 3376 3508 3384
rect 3804 3376 3812 3384
rect 3868 3376 3876 3384
rect 3996 3376 4004 3384
rect 4204 3376 4212 3384
rect 4396 3376 4404 3384
rect 4604 3376 4612 3384
rect 4684 3376 4692 3384
rect 4796 3376 4804 3384
rect 4828 3376 4836 3384
rect 4956 3376 4964 3384
rect 5004 3376 5012 3384
rect 5420 3376 5428 3384
rect 5532 3376 5540 3384
rect 5676 3376 5684 3384
rect 6060 3376 6068 3384
rect 6476 3376 6484 3384
rect 6524 3376 6532 3384
rect 6588 3376 6596 3384
rect 6668 3376 6676 3384
rect 6732 3376 6740 3384
rect 6972 3376 6980 3384
rect 7052 3376 7060 3384
rect 7196 3376 7204 3384
rect 7980 3376 7988 3384
rect 12 3356 20 3364
rect 44 3336 52 3344
rect 188 3336 196 3344
rect 252 3336 260 3344
rect 348 3336 356 3344
rect 396 3356 404 3364
rect 716 3356 724 3364
rect 444 3336 452 3344
rect 460 3336 468 3344
rect 572 3336 580 3344
rect 684 3336 692 3344
rect 700 3336 708 3344
rect 1324 3356 1332 3364
rect 1388 3356 1396 3364
rect 1756 3356 1764 3364
rect 1836 3356 1844 3364
rect 1932 3356 1940 3364
rect 2620 3356 2628 3364
rect 2636 3356 2644 3364
rect 2780 3356 2788 3364
rect 2828 3356 2836 3364
rect 2924 3356 2932 3364
rect 3420 3356 3428 3364
rect 3708 3356 3716 3364
rect 3852 3356 3860 3364
rect 3916 3356 3924 3364
rect 3932 3356 3940 3364
rect 4012 3356 4020 3364
rect 4300 3356 4308 3364
rect 4588 3356 4596 3364
rect 4780 3356 4788 3364
rect 4812 3356 4820 3364
rect 4940 3356 4948 3364
rect 5260 3356 5268 3364
rect 5452 3356 5460 3364
rect 5580 3356 5588 3364
rect 5596 3356 5604 3364
rect 5660 3356 5668 3364
rect 6396 3356 6404 3364
rect 6492 3356 6500 3364
rect 6748 3356 6756 3364
rect 7068 3356 7076 3364
rect 7084 3356 7092 3364
rect 7148 3356 7156 3364
rect 7212 3356 7220 3364
rect 7276 3356 7284 3364
rect 7500 3356 7508 3364
rect 7596 3356 7604 3364
rect 7964 3356 7972 3364
rect 8044 3356 8052 3364
rect 892 3336 900 3344
rect 988 3336 996 3344
rect 1004 3336 1012 3344
rect 1100 3336 1108 3344
rect 1532 3336 1540 3344
rect 1708 3336 1716 3344
rect 1756 3336 1764 3344
rect 1868 3336 1876 3344
rect 2012 3336 2020 3344
rect 2204 3336 2212 3344
rect 2492 3336 2500 3344
rect 2540 3336 2548 3344
rect 2556 3336 2564 3344
rect 2588 3336 2596 3344
rect 2684 3336 2692 3344
rect 2700 3336 2708 3344
rect 2796 3336 2804 3344
rect 2972 3332 2980 3340
rect 2988 3336 2996 3344
rect 3116 3336 3124 3344
rect 3164 3336 3172 3344
rect 3228 3332 3236 3340
rect 3340 3336 3348 3344
rect 3756 3336 3764 3344
rect 3788 3336 3796 3344
rect 3852 3336 3860 3344
rect 3884 3336 3892 3344
rect 3980 3336 3988 3344
rect 4028 3336 4036 3344
rect 4124 3336 4132 3344
rect 4140 3336 4148 3344
rect 4172 3336 4180 3344
rect 4236 3336 4244 3344
rect 4332 3336 4340 3344
rect 4348 3332 4356 3340
rect 4620 3336 4628 3344
rect 4716 3336 4724 3344
rect 4748 3336 4756 3344
rect 4908 3332 4916 3340
rect 5084 3336 5092 3344
rect 5148 3336 5156 3344
rect 5164 3336 5172 3344
rect 5340 3336 5348 3344
rect 5356 3336 5364 3344
rect 5404 3336 5412 3344
rect 5500 3336 5508 3344
rect 5516 3336 5524 3344
rect 5548 3336 5556 3344
rect 5804 3336 5812 3344
rect 5916 3336 5924 3344
rect 6012 3336 6020 3344
rect 6076 3336 6084 3344
rect 6108 3336 6116 3344
rect 6332 3336 6340 3344
rect 6444 3336 6452 3344
rect 6540 3336 6548 3344
rect 6556 3336 6564 3344
rect 6652 3336 6660 3344
rect 6700 3332 6708 3340
rect 6764 3336 6772 3344
rect 6892 3336 6900 3344
rect 6908 3336 6916 3344
rect 7020 3336 7028 3344
rect 7036 3336 7044 3344
rect 7644 3336 7652 3344
rect 7676 3336 7684 3344
rect 7788 3336 7796 3344
rect 7836 3336 7844 3344
rect 7852 3336 7860 3344
rect 7948 3336 7956 3344
rect 7996 3336 8004 3344
rect 8156 3336 8164 3344
rect 60 3316 68 3324
rect 92 3316 100 3324
rect 204 3316 212 3324
rect 396 3316 404 3324
rect 428 3316 436 3324
rect 524 3316 532 3324
rect 588 3316 596 3324
rect 604 3316 612 3324
rect 76 3296 84 3304
rect 140 3296 148 3304
rect 236 3296 244 3304
rect 396 3296 404 3304
rect 492 3296 500 3304
rect 508 3296 516 3304
rect 668 3316 676 3324
rect 748 3316 756 3324
rect 828 3316 836 3324
rect 892 3316 900 3324
rect 940 3316 948 3324
rect 1004 3316 1012 3324
rect 1036 3316 1044 3324
rect 1068 3316 1076 3324
rect 1132 3318 1140 3326
rect 1308 3316 1316 3324
rect 1532 3318 1540 3326
rect 1612 3316 1620 3324
rect 1676 3316 1684 3324
rect 1692 3316 1700 3324
rect 1724 3316 1732 3324
rect 1900 3316 1908 3324
rect 1980 3316 1988 3324
rect 2044 3318 2052 3326
rect 2252 3316 2260 3324
rect 2380 3316 2388 3324
rect 2460 3316 2468 3324
rect 2540 3316 2548 3324
rect 2572 3316 2580 3324
rect 2876 3316 2884 3324
rect 3068 3316 3076 3324
rect 3116 3316 3124 3324
rect 3196 3316 3204 3324
rect 3244 3316 3252 3324
rect 3260 3316 3268 3324
rect 3372 3316 3380 3324
rect 3468 3316 3476 3324
rect 3564 3318 3572 3326
rect 3628 3316 3636 3324
rect 3740 3316 3748 3324
rect 3772 3316 3780 3324
rect 3836 3316 3844 3324
rect 3916 3316 3924 3324
rect 3964 3316 3972 3324
rect 4156 3316 4164 3324
rect 4284 3316 4292 3324
rect 4460 3316 4468 3324
rect 4524 3318 4532 3326
rect 4732 3316 4740 3324
rect 4972 3316 4980 3324
rect 5036 3316 5044 3324
rect 5100 3316 5108 3324
rect 5228 3316 5236 3324
rect 5292 3316 5300 3324
rect 5324 3316 5332 3324
rect 5404 3316 5412 3324
rect 5484 3316 5492 3324
rect 5500 3316 5508 3324
rect 5564 3316 5572 3324
rect 5660 3316 5668 3324
rect 5708 3316 5716 3324
rect 636 3296 644 3304
rect 732 3296 740 3304
rect 924 3296 932 3304
rect 1068 3296 1076 3304
rect 1596 3296 1604 3304
rect 1660 3296 1668 3304
rect 1852 3296 1860 3304
rect 2428 3296 2436 3304
rect 2476 3296 2484 3304
rect 2492 3296 2500 3304
rect 2652 3296 2660 3304
rect 2748 3296 2756 3304
rect 2844 3296 2852 3304
rect 2876 3296 2884 3304
rect 3500 3296 3508 3304
rect 4060 3296 4068 3304
rect 4188 3296 4196 3304
rect 4204 3296 4212 3304
rect 76 3276 84 3284
rect 284 3276 292 3284
rect 540 3276 548 3284
rect 764 3276 772 3284
rect 780 3276 788 3284
rect 796 3276 804 3284
rect 956 3276 964 3284
rect 1628 3276 1636 3284
rect 2140 3276 2148 3284
rect 2444 3276 2452 3284
rect 3420 3276 3428 3284
rect 3708 3276 3716 3284
rect 5132 3296 5140 3304
rect 5180 3296 5188 3304
rect 5196 3296 5204 3304
rect 5388 3296 5396 3304
rect 5436 3296 5444 3304
rect 5612 3296 5620 3304
rect 5788 3316 5796 3324
rect 5884 3316 5892 3324
rect 5932 3316 5940 3324
rect 6028 3316 6036 3324
rect 6300 3318 6308 3326
rect 6108 3296 6116 3304
rect 6716 3316 6724 3324
rect 7020 3316 7028 3324
rect 7164 3316 7172 3324
rect 7356 3316 7364 3324
rect 7420 3318 7428 3326
rect 7532 3316 7540 3324
rect 7628 3316 7636 3324
rect 7692 3316 7700 3324
rect 7884 3316 7892 3324
rect 8060 3316 8068 3324
rect 8108 3316 8116 3324
rect 6364 3296 6372 3304
rect 6508 3296 6516 3304
rect 7260 3296 7268 3304
rect 7516 3296 7524 3304
rect 7596 3296 7604 3304
rect 7660 3296 7668 3304
rect 7724 3296 7732 3304
rect 7740 3296 7748 3304
rect 7772 3296 7780 3304
rect 7804 3296 7812 3304
rect 5052 3276 5060 3284
rect 5228 3276 5236 3284
rect 5740 3276 5748 3284
rect 5820 3276 5828 3284
rect 7548 3276 7556 3284
rect 7692 3276 7700 3284
rect 8092 3276 8100 3284
rect 5788 3256 5796 3264
rect 7532 3256 7540 3264
rect 12 3236 20 3244
rect 380 3236 388 3244
rect 556 3236 564 3244
rect 828 3236 836 3244
rect 1276 3236 1284 3244
rect 1356 3236 1364 3244
rect 1404 3236 1412 3244
rect 1612 3236 1620 3244
rect 2172 3236 2180 3244
rect 2364 3236 2372 3244
rect 2412 3236 2420 3244
rect 2716 3236 2724 3244
rect 4252 3236 4260 3244
rect 4316 3236 4324 3244
rect 4380 3236 4388 3244
rect 4780 3236 4788 3244
rect 5068 3236 5076 3244
rect 5100 3236 5108 3244
rect 6172 3236 6180 3244
rect 7116 3236 7124 3244
rect 7292 3236 7300 3244
rect 7484 3236 7492 3244
rect 8028 3236 8036 3244
rect 1742 3206 1750 3214
rect 1756 3206 1764 3214
rect 1770 3206 1778 3214
rect 4814 3206 4822 3214
rect 4828 3206 4836 3214
rect 4842 3206 4850 3214
rect 604 3176 612 3184
rect 732 3176 740 3184
rect 844 3176 852 3184
rect 1020 3176 1028 3184
rect 1484 3176 1492 3184
rect 1580 3176 1588 3184
rect 2492 3176 2500 3184
rect 2540 3176 2548 3184
rect 2940 3176 2948 3184
rect 4508 3176 4516 3184
rect 4556 3176 4564 3184
rect 4892 3176 4900 3184
rect 5052 3176 5060 3184
rect 5324 3176 5332 3184
rect 5500 3176 5508 3184
rect 5676 3176 5684 3184
rect 5820 3176 5828 3184
rect 5852 3176 5860 3184
rect 5900 3176 5908 3184
rect 6236 3176 6244 3184
rect 7500 3176 7508 3184
rect 7948 3176 7956 3184
rect 4460 3156 4468 3164
rect 6860 3156 6868 3164
rect 6988 3156 6996 3164
rect 60 3136 68 3144
rect 332 3136 340 3144
rect 700 3136 708 3144
rect 1228 3136 1236 3144
rect 1564 3136 1572 3144
rect 2012 3136 2020 3144
rect 2300 3136 2308 3144
rect 2412 3136 2420 3144
rect 2508 3136 2516 3144
rect 3420 3136 3428 3144
rect 3452 3136 3460 3144
rect 3580 3136 3588 3144
rect 3884 3136 3892 3144
rect 3916 3136 3924 3144
rect 4492 3136 4500 3144
rect 5100 3136 5108 3144
rect 5772 3136 5780 3144
rect 6316 3136 6324 3144
rect 6844 3136 6852 3144
rect 7036 3136 7044 3144
rect 7228 3136 7236 3144
rect 7484 3136 7492 3144
rect 7788 3136 7796 3144
rect 44 3116 52 3124
rect 316 3116 324 3124
rect 492 3116 500 3124
rect 636 3116 644 3124
rect 764 3116 772 3124
rect 1276 3116 1284 3124
rect 1340 3116 1348 3124
rect 1372 3116 1380 3124
rect 1612 3116 1620 3124
rect 1644 3116 1652 3124
rect 76 3096 84 3104
rect 92 3096 100 3104
rect 156 3096 164 3104
rect 236 3096 244 3104
rect 364 3096 372 3104
rect 732 3096 740 3104
rect 780 3096 788 3104
rect 812 3096 820 3104
rect 892 3096 900 3104
rect 1148 3096 1156 3104
rect 1164 3096 1172 3104
rect 1420 3096 1428 3104
rect 1532 3096 1540 3104
rect 1580 3096 1588 3104
rect 1660 3096 1668 3104
rect 1740 3096 1748 3104
rect 1756 3096 1764 3104
rect 1884 3116 1892 3124
rect 2076 3116 2084 3124
rect 2364 3116 2372 3124
rect 1964 3096 1972 3104
rect 2188 3096 2196 3104
rect 2364 3096 2372 3104
rect 2476 3116 2484 3124
rect 2652 3116 2660 3124
rect 2828 3116 2836 3124
rect 3196 3116 3204 3124
rect 2444 3096 2452 3104
rect 2492 3096 2500 3104
rect 2572 3096 2580 3104
rect 2636 3096 2644 3104
rect 2716 3096 2724 3104
rect 2780 3096 2788 3104
rect 3052 3096 3060 3104
rect 3148 3096 3156 3104
rect 3164 3096 3172 3104
rect 3324 3096 3332 3104
rect 3356 3096 3364 3104
rect 3452 3096 3460 3104
rect 3500 3116 3508 3124
rect 3644 3116 3652 3124
rect 3532 3096 3540 3104
rect 3564 3096 3572 3104
rect 3644 3096 3652 3104
rect 3676 3096 3684 3104
rect 3740 3116 3748 3124
rect 3852 3116 3860 3124
rect 4524 3116 4532 3124
rect 3788 3096 3796 3104
rect 3980 3096 3988 3104
rect 4300 3096 4308 3104
rect 4508 3096 4516 3104
rect 4556 3096 4564 3104
rect 4604 3116 4612 3124
rect 4668 3116 4676 3124
rect 4764 3116 4772 3124
rect 5132 3116 5140 3124
rect 5356 3116 5364 3124
rect 6172 3116 6180 3124
rect 4636 3096 4644 3104
rect 4812 3096 4820 3104
rect 4908 3096 4916 3104
rect 4956 3096 4964 3104
rect 4988 3096 4996 3104
rect 5116 3096 5124 3104
rect 5196 3094 5204 3102
rect 5532 3096 5540 3104
rect 5708 3096 5716 3104
rect 5756 3096 5764 3104
rect 5884 3096 5892 3104
rect 5932 3096 5940 3104
rect 6012 3096 6020 3104
rect 6076 3094 6084 3102
rect 6172 3096 6180 3104
rect 6204 3096 6212 3104
rect 6268 3096 6276 3104
rect 6396 3116 6404 3124
rect 6780 3116 6788 3124
rect 6876 3116 6884 3124
rect 6940 3116 6948 3124
rect 6460 3096 6468 3104
rect 6492 3096 6500 3104
rect 6508 3096 6516 3104
rect 6572 3096 6580 3104
rect 6668 3096 6676 3104
rect 6732 3096 6740 3104
rect 6860 3096 6868 3104
rect 12 3076 20 3084
rect 60 3076 68 3084
rect 108 3076 116 3084
rect 140 3076 148 3084
rect 172 3076 180 3084
rect 188 3080 196 3088
rect 60 3056 68 3064
rect 284 3076 292 3084
rect 412 3076 420 3084
rect 428 3076 436 3084
rect 524 3076 532 3084
rect 572 3076 580 3084
rect 652 3076 660 3084
rect 668 3076 676 3084
rect 716 3076 724 3084
rect 876 3076 884 3084
rect 908 3076 916 3084
rect 1052 3076 1060 3084
rect 1148 3076 1156 3084
rect 1180 3076 1188 3084
rect 1260 3076 1268 3084
rect 1276 3076 1284 3084
rect 1340 3076 1348 3084
rect 1372 3076 1380 3084
rect 1500 3076 1508 3084
rect 1612 3076 1620 3084
rect 1708 3076 1716 3084
rect 1836 3076 1844 3084
rect 1916 3076 1924 3084
rect 1980 3076 1988 3084
rect 2012 3076 2020 3084
rect 2108 3076 2116 3084
rect 2140 3076 2148 3084
rect 2460 3076 2468 3084
rect 2572 3076 2580 3084
rect 2588 3076 2596 3084
rect 2620 3076 2628 3084
rect 2684 3076 2692 3084
rect 2764 3076 2772 3084
rect 2796 3076 2804 3084
rect 2892 3076 2900 3084
rect 2924 3076 2932 3084
rect 3068 3076 3076 3084
rect 3132 3076 3140 3084
rect 3436 3076 3444 3084
rect 3548 3076 3556 3084
rect 3564 3076 3572 3084
rect 3612 3076 3620 3084
rect 3628 3076 3636 3084
rect 3676 3076 3684 3084
rect 3692 3076 3700 3084
rect 3772 3076 3780 3084
rect 3804 3076 3812 3084
rect 3836 3076 3844 3084
rect 4044 3076 4052 3084
rect 4076 3076 4084 3084
rect 4204 3076 4212 3084
rect 4236 3076 4244 3084
rect 4540 3076 4548 3084
rect 4652 3076 4660 3084
rect 4700 3076 4708 3084
rect 4716 3076 4724 3084
rect 4748 3076 4756 3084
rect 4972 3076 4980 3084
rect 5116 3076 5124 3084
rect 5564 3076 5572 3084
rect 5660 3076 5668 3084
rect 5804 3076 5812 3084
rect 5900 3076 5908 3084
rect 6108 3076 6116 3084
rect 6156 3076 6164 3084
rect 6220 3076 6228 3084
rect 6284 3076 6292 3084
rect 6300 3076 6308 3084
rect 6428 3076 6436 3084
rect 6444 3076 6452 3084
rect 6508 3076 6516 3084
rect 6684 3076 6692 3084
rect 6716 3076 6724 3084
rect 6748 3076 6756 3084
rect 6908 3096 6916 3104
rect 7084 3116 7092 3124
rect 7116 3116 7124 3124
rect 7148 3116 7156 3124
rect 7452 3116 7460 3124
rect 7516 3116 7524 3124
rect 7724 3116 7732 3124
rect 7868 3116 7876 3124
rect 7900 3116 7908 3124
rect 7932 3116 7940 3124
rect 6988 3096 6996 3104
rect 7052 3096 7060 3104
rect 7180 3096 7188 3104
rect 7292 3096 7300 3104
rect 7340 3096 7348 3104
rect 7500 3096 7508 3104
rect 7532 3096 7540 3104
rect 7596 3096 7604 3104
rect 7612 3096 7620 3104
rect 7660 3096 7668 3104
rect 7740 3096 7748 3104
rect 7804 3096 7812 3104
rect 7836 3096 7844 3104
rect 7900 3096 7908 3104
rect 8012 3096 8020 3104
rect 8028 3096 8036 3104
rect 7004 3076 7012 3084
rect 7132 3076 7140 3084
rect 7180 3076 7188 3084
rect 7356 3076 7364 3084
rect 7420 3076 7428 3084
rect 7548 3076 7556 3084
rect 7580 3076 7588 3084
rect 540 3056 548 3064
rect 620 3056 628 3064
rect 684 3056 692 3064
rect 812 3056 820 3064
rect 1212 3056 1220 3064
rect 1388 3056 1396 3064
rect 1436 3056 1444 3064
rect 1516 3056 1524 3064
rect 1820 3056 1828 3064
rect 1932 3056 1940 3064
rect 2172 3056 2180 3064
rect 2316 3056 2324 3064
rect 2556 3056 2564 3064
rect 2652 3056 2660 3064
rect 2700 3056 2708 3064
rect 2732 3056 2740 3064
rect 2908 3056 2916 3064
rect 3836 3056 3844 3064
rect 3852 3056 3860 3064
rect 4412 3056 4420 3064
rect 4428 3056 4436 3064
rect 4444 3056 4452 3064
rect 4780 3056 4788 3064
rect 4924 3056 4932 3064
rect 5068 3056 5076 3064
rect 5196 3056 5204 3064
rect 5340 3056 5348 3064
rect 5404 3056 5412 3064
rect 5420 3056 5428 3064
rect 5484 3056 5492 3064
rect 5836 3056 5844 3064
rect 6140 3056 6148 3064
rect 6588 3056 6596 3064
rect 6636 3056 6644 3064
rect 6796 3056 6804 3064
rect 7052 3056 7060 3064
rect 7756 3076 7764 3084
rect 7788 3076 7796 3084
rect 7820 3076 7828 3084
rect 7884 3076 7892 3084
rect 8028 3076 8036 3084
rect 7452 3056 7460 3064
rect 7564 3056 7572 3064
rect 7644 3056 7652 3064
rect 7676 3056 7684 3064
rect 108 3036 116 3044
rect 220 3036 228 3044
rect 252 3036 260 3044
rect 316 3036 324 3044
rect 556 3036 564 3044
rect 1196 3036 1204 3044
rect 1244 3036 1252 3044
rect 1404 3036 1412 3044
rect 1692 3036 1700 3044
rect 1804 3036 1812 3044
rect 1868 3036 1876 3044
rect 2588 3036 2596 3044
rect 2748 3036 2756 3044
rect 3868 3036 3876 3044
rect 4396 3036 4404 3044
rect 4940 3036 4948 3044
rect 5436 3036 5444 3044
rect 5612 3036 5620 3044
rect 5724 3036 5732 3044
rect 5772 3036 5780 3044
rect 5948 3036 5956 3044
rect 6556 3036 6564 3044
rect 6700 3036 6708 3044
rect 6764 3036 6772 3044
rect 6812 3036 6820 3044
rect 7628 3036 7636 3044
rect 7708 3036 7716 3044
rect 7868 3036 7876 3044
rect 7948 3036 7956 3044
rect 5340 3016 5348 3024
rect 5420 3016 5428 3024
rect 3278 3006 3286 3014
rect 3292 3006 3300 3014
rect 3306 3006 3314 3014
rect 6350 3006 6358 3014
rect 6364 3006 6372 3014
rect 6378 3006 6386 3014
rect 556 2976 564 2984
rect 764 2976 772 2984
rect 828 2976 836 2984
rect 892 2976 900 2984
rect 1324 2976 1332 2984
rect 2364 2976 2372 2984
rect 2444 2976 2452 2984
rect 3180 2976 3188 2984
rect 76 2956 84 2964
rect 92 2956 100 2964
rect 780 2956 788 2964
rect 1708 2956 1716 2964
rect 2092 2956 2100 2964
rect 2220 2956 2228 2964
rect 2492 2956 2500 2964
rect 2604 2956 2612 2964
rect 2988 2956 2996 2964
rect 3196 2956 3204 2964
rect 3436 2976 3444 2984
rect 3484 2976 3492 2984
rect 3516 2976 3524 2984
rect 3564 2976 3572 2984
rect 3596 2976 3604 2984
rect 3724 2976 3732 2984
rect 3900 2976 3908 2984
rect 4172 2976 4180 2984
rect 4972 2976 4980 2984
rect 5164 2976 5172 2984
rect 5468 2976 5476 2984
rect 5804 2976 5812 2984
rect 5996 2976 6004 2984
rect 6236 2976 6244 2984
rect 6316 2976 6324 2984
rect 6348 2976 6356 2984
rect 6636 2976 6644 2984
rect 6956 2976 6964 2984
rect 7260 2976 7268 2984
rect 7772 2976 7780 2984
rect 8060 2976 8068 2984
rect 3356 2956 3364 2964
rect 3404 2956 3412 2964
rect 3452 2956 3460 2964
rect 3532 2956 3540 2964
rect 3548 2956 3556 2964
rect 3884 2956 3892 2964
rect 4460 2956 4468 2964
rect 4588 2956 4596 2964
rect 4748 2956 4756 2964
rect 5260 2956 5268 2964
rect 5484 2956 5492 2964
rect 5660 2956 5668 2964
rect 6540 2956 6548 2964
rect 7004 2956 7012 2964
rect 7036 2956 7044 2964
rect 7116 2956 7124 2964
rect 7500 2956 7508 2964
rect 7516 2956 7524 2964
rect 7788 2956 7796 2964
rect 7932 2956 7940 2964
rect 12 2936 20 2944
rect 44 2936 52 2944
rect 188 2936 196 2944
rect 252 2936 260 2944
rect 300 2936 308 2944
rect 364 2936 372 2944
rect 588 2936 596 2944
rect 796 2936 804 2944
rect 876 2936 884 2944
rect 924 2932 932 2940
rect 940 2936 948 2944
rect 956 2936 964 2944
rect 1084 2936 1092 2944
rect 1164 2936 1172 2944
rect 1356 2936 1364 2944
rect 1388 2936 1396 2944
rect 1564 2936 1572 2944
rect 1628 2936 1636 2944
rect 1756 2936 1764 2944
rect 1804 2936 1812 2944
rect 1884 2936 1892 2944
rect 1932 2932 1940 2940
rect 2172 2936 2180 2944
rect 2300 2936 2308 2944
rect 2348 2936 2356 2944
rect 2396 2936 2404 2944
rect 2412 2932 2420 2940
rect 2556 2936 2564 2944
rect 2572 2936 2580 2944
rect 2620 2936 2628 2944
rect 2700 2936 2708 2944
rect 2796 2936 2804 2944
rect 3020 2936 3028 2944
rect 3324 2936 3332 2944
rect 3340 2936 3348 2944
rect 3372 2936 3380 2944
rect 3500 2936 3508 2944
rect 3644 2936 3652 2944
rect 3660 2936 3668 2944
rect 3756 2936 3764 2944
rect 3772 2936 3780 2944
rect 3836 2936 3844 2944
rect 3980 2936 3988 2944
rect 140 2916 148 2924
rect 156 2916 164 2924
rect 204 2916 212 2924
rect 28 2896 36 2904
rect 44 2896 52 2904
rect 172 2896 180 2904
rect 204 2896 212 2904
rect 460 2916 468 2924
rect 492 2916 500 2924
rect 636 2916 644 2924
rect 332 2896 340 2904
rect 1132 2916 1140 2924
rect 1196 2918 1204 2926
rect 1436 2916 1444 2924
rect 1580 2916 1588 2924
rect 844 2896 852 2904
rect 1660 2916 1668 2924
rect 1740 2916 1748 2924
rect 1804 2916 1812 2924
rect 1852 2916 1860 2924
rect 1884 2916 1892 2924
rect 1900 2916 1908 2924
rect 2012 2916 2020 2924
rect 2028 2916 2036 2924
rect 2044 2916 2052 2924
rect 2156 2918 2164 2926
rect 2332 2916 2340 2924
rect 2460 2916 2468 2924
rect 2508 2916 2516 2924
rect 2572 2916 2580 2924
rect 1724 2896 1732 2904
rect 2012 2896 2020 2904
rect 2380 2896 2388 2904
rect 2652 2896 2660 2904
rect 2684 2916 2692 2924
rect 2764 2918 2772 2926
rect 2924 2916 2932 2924
rect 2940 2916 2948 2924
rect 3052 2918 3060 2926
rect 3324 2916 3332 2924
rect 3580 2916 3588 2924
rect 3628 2916 3636 2924
rect 3820 2916 3828 2924
rect 3852 2916 3860 2924
rect 3932 2916 3940 2924
rect 3996 2916 4004 2924
rect 2908 2896 2916 2904
rect 3468 2896 3476 2904
rect 3804 2896 3812 2904
rect 3820 2896 3828 2904
rect 3916 2896 3924 2904
rect 3996 2896 4004 2904
rect 4076 2916 4084 2924
rect 4236 2936 4244 2944
rect 4412 2936 4420 2944
rect 4524 2936 4532 2944
rect 4556 2936 4564 2944
rect 4572 2936 4580 2944
rect 4636 2936 4644 2944
rect 4732 2936 4740 2944
rect 4124 2916 4132 2924
rect 4204 2916 4212 2924
rect 4284 2916 4292 2924
rect 4428 2916 4436 2924
rect 4044 2896 4052 2904
rect 4108 2896 4116 2904
rect 4508 2916 4516 2924
rect 4620 2916 4628 2924
rect 4684 2916 4692 2924
rect 4796 2916 4804 2924
rect 4860 2936 4868 2944
rect 4956 2936 4964 2944
rect 5020 2936 5028 2944
rect 5164 2936 5172 2944
rect 5308 2936 5316 2944
rect 5532 2936 5540 2944
rect 5548 2936 5556 2944
rect 5708 2936 5716 2944
rect 5788 2936 5796 2944
rect 5916 2936 5924 2944
rect 6108 2936 6116 2944
rect 6188 2936 6196 2944
rect 6508 2936 6516 2944
rect 6620 2936 6628 2944
rect 6748 2936 6756 2944
rect 6828 2936 6836 2944
rect 6940 2936 6948 2944
rect 6988 2936 6996 2944
rect 7036 2936 7044 2944
rect 7084 2936 7092 2944
rect 7132 2936 7140 2944
rect 7228 2936 7236 2944
rect 7372 2936 7380 2944
rect 7388 2936 7396 2944
rect 7436 2936 7444 2944
rect 7548 2936 7556 2944
rect 7660 2936 7668 2944
rect 7724 2936 7732 2944
rect 5004 2916 5012 2924
rect 5068 2916 5076 2924
rect 5148 2916 5156 2924
rect 5356 2916 5364 2924
rect 5516 2916 5524 2924
rect 5612 2916 5620 2924
rect 5708 2916 5716 2924
rect 5756 2916 5764 2924
rect 5900 2916 5908 2924
rect 6092 2916 6100 2924
rect 6204 2916 6212 2924
rect 6252 2916 6260 2924
rect 6476 2918 6484 2926
rect 6572 2916 6580 2924
rect 6588 2916 6596 2924
rect 6604 2916 6612 2924
rect 6764 2918 6772 2926
rect 6844 2916 6852 2924
rect 6860 2916 6868 2924
rect 4476 2896 4484 2904
rect 4540 2896 4548 2904
rect 4604 2896 4612 2904
rect 4700 2896 4708 2904
rect 5580 2896 5588 2904
rect 5724 2896 5732 2904
rect 5740 2896 5748 2904
rect 6572 2896 6580 2904
rect 6924 2916 6932 2924
rect 7036 2916 7044 2924
rect 7068 2916 7076 2924
rect 7132 2916 7140 2924
rect 7404 2916 7412 2924
rect 6892 2896 6900 2904
rect 6956 2896 6964 2904
rect 7452 2916 7460 2924
rect 7468 2916 7476 2924
rect 7596 2916 7604 2924
rect 7628 2916 7636 2924
rect 7740 2916 7748 2924
rect 7836 2916 7844 2924
rect 7932 2918 7940 2926
rect 8076 2916 8084 2924
rect 7484 2896 7492 2904
rect 7836 2896 7844 2904
rect 7868 2896 7876 2904
rect 236 2876 244 2884
rect 748 2876 756 2884
rect 1292 2876 1300 2884
rect 1548 2876 1556 2884
rect 1612 2876 1620 2884
rect 1948 2876 1956 2884
rect 2524 2876 2532 2884
rect 2892 2876 2900 2884
rect 3948 2876 3956 2884
rect 4140 2876 4148 2884
rect 4364 2876 4372 2884
rect 4396 2876 4404 2884
rect 5020 2876 5028 2884
rect 5212 2876 5220 2884
rect 5692 2876 5700 2884
rect 5740 2876 5748 2884
rect 6668 2876 6676 2884
rect 7516 2876 7524 2884
rect 8156 2876 8164 2884
rect 3420 2856 3428 2864
rect 268 2836 276 2844
rect 1100 2836 1108 2844
rect 2284 2836 2292 2844
rect 2300 2836 2308 2844
rect 3964 2836 3972 2844
rect 4124 2836 4132 2844
rect 4668 2836 4676 2844
rect 4748 2836 4756 2844
rect 5100 2836 5108 2844
rect 5276 2836 5284 2844
rect 5500 2836 5508 2844
rect 5644 2836 5652 2844
rect 6236 2836 6244 2844
rect 7116 2836 7124 2844
rect 1742 2806 1750 2814
rect 1756 2806 1764 2814
rect 1770 2806 1778 2814
rect 4814 2806 4822 2814
rect 4828 2806 4836 2814
rect 4842 2806 4850 2814
rect 188 2776 196 2784
rect 204 2776 212 2784
rect 732 2776 740 2784
rect 828 2776 836 2784
rect 844 2776 852 2784
rect 1548 2776 1556 2784
rect 2668 2776 2676 2784
rect 2860 2776 2868 2784
rect 2876 2776 2884 2784
rect 2924 2776 2932 2784
rect 3244 2776 3252 2784
rect 4092 2776 4100 2784
rect 4572 2776 4580 2784
rect 5756 2776 5764 2784
rect 5820 2776 5828 2784
rect 6972 2776 6980 2784
rect 6988 2776 6996 2784
rect 7884 2776 7892 2784
rect 7932 2776 7940 2784
rect 1884 2756 1892 2764
rect 4764 2756 4772 2764
rect 7420 2756 7428 2764
rect 748 2736 756 2744
rect 892 2736 900 2744
rect 1388 2736 1396 2744
rect 1420 2736 1428 2744
rect 4060 2736 4068 2744
rect 4684 2736 4692 2744
rect 4796 2736 4804 2744
rect 4892 2736 4900 2744
rect 5516 2736 5524 2744
rect 5692 2736 5700 2744
rect 6108 2736 6116 2744
rect 6172 2736 6180 2744
rect 6204 2736 6212 2744
rect 7964 2736 7972 2744
rect 8092 2736 8100 2744
rect 396 2716 404 2724
rect 428 2716 436 2724
rect 1116 2716 1124 2724
rect 1164 2716 1172 2724
rect 1580 2716 1588 2724
rect 1612 2716 1620 2724
rect 1644 2716 1652 2724
rect 1772 2716 1780 2724
rect 1868 2716 1876 2724
rect 3196 2716 3204 2724
rect 3548 2716 3556 2724
rect 3724 2716 3732 2724
rect 60 2694 68 2702
rect 124 2696 132 2704
rect 268 2696 276 2704
rect 316 2696 324 2704
rect 428 2696 436 2704
rect 508 2696 516 2704
rect 604 2694 612 2702
rect 828 2696 836 2704
rect 876 2696 884 2704
rect 892 2696 900 2704
rect 1068 2696 1076 2704
rect 1308 2696 1316 2704
rect 1612 2696 1620 2704
rect 1628 2696 1636 2704
rect 1692 2696 1700 2704
rect 1820 2696 1828 2704
rect 1916 2696 1924 2704
rect 2044 2696 2052 2704
rect 2076 2696 2084 2704
rect 2092 2696 2100 2704
rect 2172 2696 2180 2704
rect 2364 2696 2372 2704
rect 2476 2696 2484 2704
rect 2668 2696 2676 2704
rect 2732 2694 2740 2702
rect 2908 2696 2916 2704
rect 2988 2696 2996 2704
rect 3052 2694 3060 2702
rect 3164 2696 3172 2704
rect 3180 2696 3188 2704
rect 3388 2694 3396 2702
rect 3452 2696 3460 2704
rect 3580 2696 3588 2704
rect 3708 2696 3716 2704
rect 3836 2716 3844 2724
rect 4268 2716 4276 2724
rect 4316 2716 4324 2724
rect 3964 2696 3972 2704
rect 4236 2696 4244 2704
rect 4540 2716 4548 2724
rect 5164 2716 5172 2724
rect 5324 2716 5332 2724
rect 5468 2716 5476 2724
rect 5484 2716 5492 2724
rect 5644 2716 5652 2724
rect 4412 2696 4420 2704
rect 4444 2696 4452 2704
rect 4492 2696 4500 2704
rect 4556 2696 4564 2704
rect 4620 2696 4628 2704
rect 4668 2696 4676 2704
rect 4716 2696 4724 2704
rect 4748 2696 4756 2704
rect 4956 2696 4964 2704
rect 5004 2696 5012 2704
rect 5132 2696 5140 2704
rect 5148 2696 5156 2704
rect 5180 2696 5188 2704
rect 5244 2696 5252 2704
rect 5292 2696 5300 2704
rect 5308 2696 5316 2704
rect 5564 2696 5572 2704
rect 5596 2696 5604 2704
rect 5852 2716 5860 2724
rect 5692 2696 5700 2704
rect 5772 2696 5780 2704
rect 5820 2696 5828 2704
rect 5868 2696 5876 2704
rect 5900 2696 5908 2704
rect 5932 2696 5940 2704
rect 5948 2696 5956 2704
rect 6044 2696 6052 2704
rect 7212 2716 7220 2724
rect 6140 2696 6148 2704
rect 6268 2696 6276 2704
rect 6636 2696 6644 2704
rect 6732 2696 6740 2704
rect 6940 2696 6948 2704
rect 7052 2696 7060 2704
rect 7564 2716 7572 2724
rect 7804 2716 7812 2724
rect 7868 2716 7876 2724
rect 7996 2716 8004 2724
rect 8012 2716 8020 2724
rect 8060 2716 8068 2724
rect 7116 2694 7124 2702
rect 7260 2696 7268 2704
rect 7324 2696 7332 2704
rect 7356 2696 7364 2704
rect 7388 2696 7396 2704
rect 7404 2696 7412 2704
rect 7468 2696 7476 2704
rect 7484 2696 7492 2704
rect 7516 2696 7524 2704
rect 7548 2696 7556 2704
rect 7676 2696 7684 2704
rect 7804 2696 7812 2704
rect 7836 2696 7844 2704
rect 7964 2696 7972 2704
rect 28 2676 36 2684
rect 476 2676 484 2684
rect 572 2676 580 2684
rect 780 2676 788 2684
rect 924 2676 932 2684
rect 1052 2676 1060 2684
rect 1084 2676 1092 2684
rect 1132 2676 1140 2684
rect 1228 2676 1236 2684
rect 1292 2676 1300 2684
rect 1404 2676 1412 2684
rect 1436 2676 1444 2684
rect 1628 2676 1636 2684
rect 1836 2676 1844 2684
rect 1948 2676 1956 2684
rect 2012 2676 2020 2684
rect 2060 2676 2068 2684
rect 2124 2676 2132 2684
rect 2140 2676 2148 2684
rect 2236 2676 2244 2684
rect 2412 2676 2420 2684
rect 2492 2676 2500 2684
rect 2620 2676 2628 2684
rect 2700 2676 2708 2684
rect 2796 2676 2804 2684
rect 3020 2676 3028 2684
rect 3372 2676 3380 2684
rect 3484 2676 3492 2684
rect 3500 2676 3508 2684
rect 3596 2676 3604 2684
rect 3692 2676 3700 2684
rect 3724 2676 3732 2684
rect 3756 2676 3764 2684
rect 3788 2676 3796 2684
rect 3868 2676 3876 2684
rect 3900 2676 3908 2684
rect 4076 2676 4084 2684
rect 4204 2676 4212 2684
rect 4220 2676 4228 2684
rect 4284 2676 4292 2684
rect 4364 2676 4372 2684
rect 4380 2676 4388 2684
rect 4508 2676 4516 2684
rect 4556 2676 4564 2684
rect 4732 2676 4740 2684
rect 4828 2676 4836 2684
rect 5180 2676 5188 2684
rect 5212 2676 5220 2684
rect 5228 2676 5236 2684
rect 5356 2676 5364 2684
rect 5388 2676 5396 2684
rect 5436 2676 5444 2684
rect 5516 2676 5524 2684
rect 5580 2676 5588 2684
rect 5596 2676 5604 2684
rect 5708 2676 5716 2684
rect 5884 2676 5892 2684
rect 5916 2676 5924 2684
rect 5980 2680 5988 2688
rect 5996 2676 6004 2684
rect 6092 2676 6100 2684
rect 6156 2676 6164 2684
rect 6332 2676 6340 2684
rect 6412 2676 6420 2684
rect 6508 2676 6516 2684
rect 6684 2676 6692 2684
rect 6716 2676 6724 2684
rect 6780 2676 6788 2684
rect 6908 2676 6916 2684
rect 6924 2676 6932 2684
rect 7068 2676 7076 2684
rect 7180 2676 7188 2684
rect 7340 2676 7348 2684
rect 7372 2676 7380 2684
rect 7420 2676 7428 2684
rect 7452 2676 7460 2684
rect 7484 2676 7492 2684
rect 7532 2676 7540 2684
rect 7580 2676 7588 2684
rect 7596 2676 7604 2684
rect 7660 2676 7668 2684
rect 7852 2676 7860 2684
rect 7900 2676 7908 2684
rect 7948 2676 7956 2684
rect 8044 2676 8052 2684
rect 8092 2676 8100 2684
rect 476 2656 484 2664
rect 764 2656 772 2664
rect 796 2656 804 2664
rect 940 2656 948 2664
rect 1004 2656 1012 2664
rect 1020 2656 1028 2664
rect 1724 2656 1732 2664
rect 1788 2656 1796 2664
rect 1980 2656 1988 2664
rect 2028 2656 2036 2664
rect 2636 2656 2644 2664
rect 3116 2656 3124 2664
rect 3452 2656 3460 2664
rect 3532 2656 3540 2664
rect 4460 2656 4468 2664
rect 4556 2656 4564 2664
rect 4588 2656 4596 2664
rect 4636 2656 4644 2664
rect 4652 2656 4660 2664
rect 5084 2656 5092 2664
rect 5260 2656 5268 2664
rect 5724 2656 5732 2664
rect 5756 2656 5764 2664
rect 6012 2656 6020 2664
rect 7308 2656 7316 2664
rect 7916 2656 7924 2664
rect 8124 2656 8132 2664
rect 540 2636 548 2644
rect 732 2636 740 2644
rect 956 2636 964 2644
rect 1036 2636 1044 2644
rect 1100 2636 1108 2644
rect 1964 2636 1972 2644
rect 2252 2636 2260 2644
rect 2444 2636 2452 2644
rect 2876 2636 2884 2644
rect 3564 2636 3572 2644
rect 4268 2636 4276 2644
rect 4604 2636 4612 2644
rect 4764 2636 4772 2644
rect 5484 2636 5492 2644
rect 6444 2636 6452 2644
rect 6524 2636 6532 2644
rect 6764 2636 6772 2644
rect 6972 2636 6980 2644
rect 7228 2636 7236 2644
rect 8012 2636 8020 2644
rect 8108 2636 8116 2644
rect 940 2616 948 2624
rect 3278 2606 3286 2614
rect 3292 2606 3300 2614
rect 3306 2606 3314 2614
rect 6350 2606 6358 2614
rect 6364 2606 6372 2614
rect 6378 2606 6386 2614
rect 1996 2596 2004 2604
rect 2652 2596 2660 2604
rect 28 2576 36 2584
rect 844 2576 852 2584
rect 1500 2576 1508 2584
rect 1980 2576 1988 2584
rect 2380 2576 2388 2584
rect 2524 2576 2532 2584
rect 2556 2576 2564 2584
rect 2956 2576 2964 2584
rect 3196 2576 3204 2584
rect 3452 2576 3460 2584
rect 3788 2576 3796 2584
rect 3836 2576 3844 2584
rect 4140 2576 4148 2584
rect 4172 2576 4180 2584
rect 4476 2576 4484 2584
rect 4620 2576 4628 2584
rect 5116 2576 5124 2584
rect 5164 2576 5172 2584
rect 5180 2576 5188 2584
rect 5228 2576 5236 2584
rect 5548 2576 5556 2584
rect 5708 2576 5716 2584
rect 5772 2576 5780 2584
rect 6044 2576 6052 2584
rect 6428 2576 6436 2584
rect 6652 2576 6660 2584
rect 6940 2576 6948 2584
rect 6956 2576 6964 2584
rect 7468 2576 7476 2584
rect 7580 2576 7588 2584
rect 8108 2576 8116 2584
rect 540 2556 548 2564
rect 780 2556 788 2564
rect 924 2556 932 2564
rect 1004 2556 1012 2564
rect 1228 2556 1236 2564
rect 1388 2556 1396 2564
rect 1484 2556 1492 2564
rect 1516 2556 1524 2564
rect 1996 2556 2004 2564
rect 2060 2556 2068 2564
rect 2220 2556 2228 2564
rect 2460 2556 2468 2564
rect 2572 2556 2580 2564
rect 2588 2556 2596 2564
rect 2652 2556 2660 2564
rect 2796 2556 2804 2564
rect 3100 2556 3108 2564
rect 3116 2556 3124 2564
rect 3148 2556 3156 2564
rect 3420 2556 3428 2564
rect 3468 2556 3476 2564
rect 3820 2556 3828 2564
rect 3964 2556 3972 2564
rect 4028 2556 4036 2564
rect 4156 2556 4164 2564
rect 4300 2556 4308 2564
rect 4428 2556 4436 2564
rect 4556 2556 4564 2564
rect 4572 2556 4580 2564
rect 4748 2556 4756 2564
rect 140 2536 148 2544
rect 268 2536 276 2544
rect 508 2536 516 2544
rect 620 2536 628 2544
rect 796 2536 804 2544
rect 892 2536 900 2544
rect 988 2536 996 2544
rect 1084 2536 1092 2544
rect 1100 2536 1108 2544
rect 1148 2536 1156 2544
rect 1308 2536 1316 2544
rect 1340 2536 1348 2544
rect 1452 2536 1460 2544
rect 1564 2536 1572 2544
rect 1596 2536 1604 2544
rect 1676 2536 1684 2544
rect 1692 2536 1700 2544
rect 1740 2536 1748 2544
rect 1932 2536 1940 2544
rect 2076 2536 2084 2544
rect 2364 2536 2372 2544
rect 2476 2536 2484 2544
rect 2860 2536 2868 2544
rect 2908 2536 2916 2544
rect 2972 2536 2980 2544
rect 3020 2536 3028 2544
rect 3084 2536 3092 2544
rect 3180 2536 3188 2544
rect 3212 2536 3220 2544
rect 3308 2536 3316 2544
rect 3388 2536 3396 2544
rect 3484 2536 3492 2544
rect 3596 2536 3604 2544
rect 3804 2536 3812 2544
rect 3868 2532 3876 2540
rect 3884 2536 3892 2544
rect 4092 2536 4100 2544
rect 4204 2536 4212 2544
rect 4396 2536 4404 2544
rect 4444 2536 4452 2544
rect 4588 2536 4596 2544
rect 4636 2536 4644 2544
rect 4684 2536 4692 2544
rect 5132 2536 5140 2544
rect 5324 2556 5332 2564
rect 5404 2556 5412 2564
rect 5580 2556 5588 2564
rect 5660 2556 5668 2564
rect 5724 2556 5732 2564
rect 5212 2536 5220 2544
rect 5260 2536 5268 2544
rect 5500 2536 5508 2544
rect 5516 2536 5524 2544
rect 5564 2536 5572 2544
rect 5644 2536 5652 2544
rect 5756 2536 5764 2544
rect 5868 2556 5876 2564
rect 6140 2556 6148 2564
rect 6156 2556 6164 2564
rect 6236 2556 6244 2564
rect 6748 2556 6756 2564
rect 7276 2556 7284 2564
rect 7596 2556 7604 2564
rect 7612 2556 7620 2564
rect 7644 2556 7652 2564
rect 7676 2556 7684 2564
rect 7740 2556 7748 2564
rect 7916 2556 7924 2564
rect 5852 2536 5860 2544
rect 5964 2536 5972 2544
rect 6028 2536 6036 2544
rect 6124 2536 6132 2544
rect 6204 2536 6212 2544
rect 6252 2536 6260 2544
rect 6348 2536 6356 2544
rect 6588 2536 6596 2544
rect 6780 2536 6788 2544
rect 7116 2536 7124 2544
rect 7148 2536 7156 2544
rect 7356 2536 7364 2544
rect 7564 2536 7572 2544
rect 284 2518 292 2526
rect 476 2518 484 2526
rect 604 2516 612 2524
rect 812 2516 820 2524
rect 844 2516 852 2524
rect 892 2516 900 2524
rect 1068 2516 1076 2524
rect 1100 2516 1108 2524
rect 1164 2516 1172 2524
rect 1180 2516 1188 2524
rect 1260 2516 1268 2524
rect 1356 2516 1364 2524
rect 1404 2516 1412 2524
rect 1468 2516 1476 2524
rect 1548 2516 1556 2524
rect 1612 2516 1620 2524
rect 1660 2516 1668 2524
rect 1724 2516 1732 2524
rect 1836 2516 1844 2524
rect 1900 2516 1908 2524
rect 1948 2516 1956 2524
rect 1980 2516 1988 2524
rect 2252 2516 2260 2524
rect 2348 2516 2356 2524
rect 2428 2516 2436 2524
rect 2492 2516 2500 2524
rect 2540 2516 2548 2524
rect 2796 2518 2804 2526
rect 2988 2516 2996 2524
rect 844 2496 852 2504
rect 860 2496 868 2504
rect 924 2496 932 2504
rect 972 2496 980 2504
rect 1020 2496 1028 2504
rect 1036 2496 1044 2504
rect 1260 2496 1268 2504
rect 1340 2496 1348 2504
rect 1628 2496 1636 2504
rect 1692 2496 1700 2504
rect 1852 2496 1860 2504
rect 1916 2496 1924 2504
rect 2364 2496 2372 2504
rect 2892 2496 2900 2504
rect 2956 2496 2964 2504
rect 3132 2516 3140 2524
rect 3164 2516 3172 2524
rect 3228 2516 3236 2524
rect 3260 2516 3268 2524
rect 3436 2516 3444 2524
rect 3500 2516 3508 2524
rect 3036 2496 3044 2504
rect 3244 2496 3252 2504
rect 3356 2496 3364 2504
rect 3420 2496 3428 2504
rect 3532 2496 3540 2504
rect 3580 2516 3588 2524
rect 3660 2518 3668 2526
rect 3708 2516 3716 2524
rect 4012 2516 4020 2524
rect 4108 2516 4116 2524
rect 4188 2516 4196 2524
rect 4252 2516 4260 2524
rect 4268 2516 4276 2524
rect 4348 2496 4356 2504
rect 4380 2516 4388 2524
rect 4524 2516 4532 2524
rect 4652 2516 4660 2524
rect 4748 2518 4756 2526
rect 5004 2516 5012 2524
rect 5036 2516 5044 2524
rect 4476 2496 4484 2504
rect 4540 2496 4548 2504
rect 4684 2496 4692 2504
rect 5276 2516 5284 2524
rect 5308 2496 5316 2504
rect 5356 2516 5364 2524
rect 5452 2516 5460 2524
rect 5564 2496 5572 2504
rect 5692 2516 5700 2524
rect 5740 2516 5748 2524
rect 5804 2516 5812 2524
rect 5852 2516 5860 2524
rect 5932 2516 5940 2524
rect 5980 2516 5988 2524
rect 6028 2516 6036 2524
rect 6108 2516 6116 2524
rect 6252 2516 6260 2524
rect 6268 2516 6276 2524
rect 6300 2516 6308 2524
rect 6364 2516 6372 2524
rect 6540 2516 6548 2524
rect 6620 2516 6628 2524
rect 6684 2516 6692 2524
rect 6700 2516 6708 2524
rect 6812 2518 6820 2526
rect 7084 2518 7092 2526
rect 5612 2496 5620 2504
rect 5884 2496 5892 2504
rect 5948 2496 5956 2504
rect 6012 2496 6020 2504
rect 6060 2496 6068 2504
rect 6076 2496 6084 2504
rect 6172 2496 6180 2504
rect 6204 2496 6212 2504
rect 6300 2496 6308 2504
rect 6668 2496 6676 2504
rect 7180 2496 7188 2504
rect 7212 2516 7220 2524
rect 7244 2516 7252 2524
rect 7340 2518 7348 2526
rect 7788 2536 7796 2544
rect 7804 2536 7812 2544
rect 7884 2536 7892 2544
rect 7500 2516 7508 2524
rect 7548 2516 7556 2524
rect 7628 2516 7636 2524
rect 7676 2516 7684 2524
rect 7708 2516 7716 2524
rect 7740 2516 7748 2524
rect 7820 2516 7828 2524
rect 8012 2516 8020 2524
rect 8028 2516 8036 2524
rect 7484 2496 7492 2504
rect 7740 2496 7748 2504
rect 7756 2496 7764 2504
rect 7804 2496 7812 2504
rect 1532 2476 1540 2484
rect 1820 2476 1828 2484
rect 1884 2476 1892 2484
rect 3276 2476 3284 2484
rect 3580 2476 3588 2484
rect 4396 2476 4404 2484
rect 4508 2476 4516 2484
rect 4524 2476 4532 2484
rect 4556 2476 4564 2484
rect 4620 2476 4628 2484
rect 5404 2476 5412 2484
rect 5916 2476 5924 2484
rect 7516 2476 7524 2484
rect 1660 2456 1668 2464
rect 1836 2456 1844 2464
rect 6220 2456 6228 2464
rect 28 2436 36 2444
rect 156 2436 164 2444
rect 348 2436 356 2444
rect 556 2436 564 2444
rect 572 2436 580 2444
rect 732 2436 740 2444
rect 1068 2436 1076 2444
rect 1116 2436 1124 2444
rect 1420 2436 1428 2444
rect 1564 2436 1572 2444
rect 1900 2436 1908 2444
rect 2188 2436 2196 2444
rect 2284 2436 2292 2444
rect 2636 2436 2644 2444
rect 2668 2436 2676 2444
rect 3260 2436 3268 2444
rect 3900 2436 3908 2444
rect 4236 2436 4244 2444
rect 4524 2436 4532 2444
rect 4876 2436 4884 2444
rect 5932 2436 5940 2444
rect 6108 2436 6116 2444
rect 6652 2436 6660 2444
rect 7500 2436 7508 2444
rect 7916 2436 7924 2444
rect 1742 2406 1750 2414
rect 1756 2406 1764 2414
rect 1770 2406 1778 2414
rect 4814 2406 4822 2414
rect 4828 2406 4836 2414
rect 4842 2406 4850 2414
rect 300 2376 308 2384
rect 844 2376 852 2384
rect 2124 2376 2132 2384
rect 2684 2376 2692 2384
rect 2876 2376 2884 2384
rect 3052 2376 3060 2384
rect 3196 2376 3204 2384
rect 3532 2376 3540 2384
rect 3692 2376 3700 2384
rect 3932 2376 3940 2384
rect 4140 2376 4148 2384
rect 5212 2376 5220 2384
rect 6300 2376 6308 2384
rect 6700 2376 6708 2384
rect 7468 2376 7476 2384
rect 7900 2376 7908 2384
rect 364 2356 372 2364
rect 508 2356 516 2364
rect 1052 2356 1060 2364
rect 3916 2356 3924 2364
rect 5836 2356 5844 2364
rect 6668 2356 6676 2364
rect 7340 2356 7348 2364
rect 316 2336 324 2344
rect 380 2336 388 2344
rect 652 2336 660 2344
rect 1068 2336 1076 2344
rect 1116 2336 1124 2344
rect 1516 2336 1524 2344
rect 2844 2336 2852 2344
rect 2892 2336 2900 2344
rect 3276 2336 3284 2344
rect 4508 2336 4516 2344
rect 4588 2336 4596 2344
rect 5820 2336 5828 2344
rect 268 2316 276 2324
rect 284 2316 292 2324
rect 348 2316 356 2324
rect 444 2316 452 2324
rect 540 2316 548 2324
rect 604 2316 612 2324
rect 1036 2316 1044 2324
rect 1148 2316 1156 2324
rect 1212 2316 1220 2324
rect 1228 2316 1236 2324
rect 1260 2316 1268 2324
rect 1436 2316 1444 2324
rect 1532 2316 1540 2324
rect 2060 2316 2068 2324
rect 2620 2316 2628 2324
rect 2732 2316 2740 2324
rect 2796 2316 2804 2324
rect 76 2296 84 2304
rect 300 2296 308 2304
rect 364 2296 372 2304
rect 508 2296 516 2304
rect 540 2296 548 2304
rect 604 2296 612 2304
rect 732 2296 740 2304
rect 764 2296 772 2304
rect 972 2294 980 2302
rect 1052 2296 1060 2304
rect 1100 2296 1108 2304
rect 1132 2296 1140 2304
rect 1180 2296 1188 2304
rect 1308 2296 1316 2304
rect 1356 2296 1364 2304
rect 1388 2296 1396 2304
rect 1548 2296 1556 2304
rect 1564 2296 1572 2304
rect 1692 2296 1700 2304
rect 1868 2296 1876 2304
rect 1900 2296 1908 2304
rect 1948 2296 1956 2304
rect 2028 2296 2036 2304
rect 2060 2296 2068 2304
rect 2188 2296 2196 2304
rect 2236 2296 2244 2304
rect 2460 2296 2468 2304
rect 2636 2296 2644 2304
rect 2716 2296 2724 2304
rect 2764 2296 2772 2304
rect 2924 2316 2932 2324
rect 3004 2316 3012 2324
rect 3244 2316 3252 2324
rect 3980 2316 3988 2324
rect 4332 2316 4340 2324
rect 4412 2316 4420 2324
rect 4556 2316 4564 2324
rect 4636 2316 4644 2324
rect 4700 2316 4708 2324
rect 2844 2296 2852 2304
rect 2908 2296 2916 2304
rect 3100 2296 3108 2304
rect 3148 2296 3156 2304
rect 3228 2296 3236 2304
rect 3260 2296 3268 2304
rect 3340 2296 3348 2304
rect 3404 2294 3412 2302
rect 3468 2296 3476 2304
rect 3548 2296 3556 2304
rect 3724 2296 3732 2304
rect 3804 2296 3812 2304
rect 3964 2296 3972 2304
rect 3996 2296 4004 2304
rect 4012 2296 4020 2304
rect 4092 2296 4100 2304
rect 4268 2294 4276 2302
rect 4364 2296 4372 2304
rect 4396 2296 4404 2304
rect 4460 2296 4468 2304
rect 4572 2296 4580 2304
rect 4668 2296 4676 2304
rect 4780 2316 4788 2324
rect 4844 2316 4852 2324
rect 5020 2316 5028 2324
rect 5068 2316 5076 2324
rect 5436 2316 5444 2324
rect 5500 2316 5508 2324
rect 5612 2316 5620 2324
rect 4748 2296 4756 2304
rect 4812 2296 4820 2304
rect 4924 2296 4932 2304
rect 5004 2296 5012 2304
rect 5084 2296 5092 2304
rect 5244 2296 5252 2304
rect 5628 2296 5636 2304
rect 5644 2296 5652 2304
rect 5676 2296 5684 2304
rect 5740 2296 5748 2304
rect 5756 2296 5764 2304
rect 5820 2296 5828 2304
rect 5916 2336 5924 2344
rect 6092 2336 6100 2344
rect 6284 2336 6292 2344
rect 7228 2336 7236 2344
rect 7804 2336 7812 2344
rect 7884 2336 7892 2344
rect 8108 2336 8116 2344
rect 5852 2316 5860 2324
rect 6060 2316 6068 2324
rect 6124 2316 6132 2324
rect 6204 2316 6212 2324
rect 6316 2316 6324 2324
rect 6428 2316 6436 2324
rect 6796 2316 6804 2324
rect 6812 2316 6820 2324
rect 6860 2316 6868 2324
rect 6876 2316 6884 2324
rect 6940 2316 6948 2324
rect 6012 2296 6020 2304
rect 6076 2296 6084 2304
rect 6124 2296 6132 2304
rect 6156 2296 6164 2304
rect 6300 2296 6308 2304
rect 6540 2294 6548 2302
rect 6588 2296 6596 2304
rect 6684 2296 6692 2304
rect 6748 2296 6756 2304
rect 6988 2316 6996 2324
rect 7244 2316 7252 2324
rect 7500 2316 7508 2324
rect 7564 2316 7572 2324
rect 7596 2316 7604 2324
rect 7692 2316 7700 2324
rect 6988 2296 6996 2304
rect 7116 2296 7124 2304
rect 7372 2296 7380 2304
rect 7404 2296 7412 2304
rect 7468 2296 7476 2304
rect 7500 2296 7508 2304
rect 7548 2296 7556 2304
rect 7660 2296 7668 2304
rect 7772 2316 7780 2324
rect 7724 2296 7732 2304
rect 7740 2296 7748 2304
rect 7788 2296 7796 2304
rect 7980 2294 7988 2302
rect 8028 2296 8036 2304
rect 28 2276 36 2284
rect 236 2276 244 2284
rect 412 2276 420 2284
rect 556 2276 564 2284
rect 812 2276 820 2284
rect 940 2276 948 2284
rect 1004 2276 1012 2284
rect 1164 2276 1172 2284
rect 1196 2276 1204 2284
rect 1292 2276 1300 2284
rect 1404 2276 1412 2284
rect 1468 2276 1476 2284
rect 1644 2276 1652 2284
rect 1964 2276 1972 2284
rect 2412 2276 2420 2284
rect 2588 2276 2596 2284
rect 2652 2276 2660 2284
rect 2684 2276 2692 2284
rect 2748 2276 2756 2284
rect 2860 2276 2868 2284
rect 2956 2276 2964 2284
rect 2988 2276 2996 2284
rect 3036 2276 3044 2284
rect 3084 2276 3092 2284
rect 3340 2276 3348 2284
rect 3372 2276 3380 2284
rect 3676 2276 3684 2284
rect 3756 2276 3764 2284
rect 4076 2276 4084 2284
rect 4236 2276 4244 2284
rect 4380 2276 4388 2284
rect 4412 2276 4420 2284
rect 4444 2276 4452 2284
rect 4540 2276 4548 2284
rect 4652 2276 4660 2284
rect 4716 2276 4724 2284
rect 4764 2276 4772 2284
rect 4828 2276 4836 2284
rect 4940 2276 4948 2284
rect 4988 2276 4996 2284
rect 5052 2276 5060 2284
rect 5260 2276 5268 2284
rect 5404 2276 5412 2284
rect 5452 2276 5460 2284
rect 5484 2276 5492 2284
rect 5516 2276 5524 2284
rect 5580 2280 5588 2288
rect 5596 2276 5604 2284
rect 5660 2276 5668 2284
rect 5692 2276 5700 2284
rect 5724 2276 5732 2284
rect 5788 2276 5796 2284
rect 5900 2276 5908 2284
rect 6028 2276 6036 2284
rect 6172 2276 6180 2284
rect 6700 2276 6708 2284
rect 6732 2276 6740 2284
rect 6764 2276 6772 2284
rect 6860 2276 6868 2284
rect 6892 2276 6900 2284
rect 6908 2276 6916 2284
rect 7068 2276 7076 2284
rect 7164 2276 7172 2284
rect 7276 2276 7284 2284
rect 7356 2276 7364 2284
rect 220 2256 228 2264
rect 476 2256 484 2264
rect 636 2256 644 2264
rect 1244 2256 1252 2264
rect 1340 2256 1348 2264
rect 1612 2256 1620 2264
rect 1820 2256 1828 2264
rect 1900 2256 1908 2264
rect 1980 2256 1988 2264
rect 2108 2256 2116 2264
rect 2316 2256 2324 2264
rect 2380 2256 2388 2264
rect 2716 2256 2724 2264
rect 3052 2256 3060 2264
rect 3164 2256 3172 2264
rect 4060 2256 4068 2264
rect 4476 2256 4484 2264
rect 4620 2256 4628 2264
rect 4780 2256 4788 2264
rect 4956 2256 4964 2264
rect 5020 2256 5028 2264
rect 5084 2256 5092 2264
rect 5532 2256 5540 2264
rect 5884 2256 5892 2264
rect 5964 2256 5972 2264
rect 6188 2256 6196 2264
rect 6252 2256 6260 2264
rect 6332 2256 6340 2264
rect 6444 2256 6452 2264
rect 6460 2256 6468 2264
rect 7036 2256 7044 2264
rect 7292 2256 7300 2264
rect 7356 2256 7364 2264
rect 7452 2276 7460 2284
rect 7644 2276 7652 2284
rect 7756 2276 7764 2284
rect 7852 2276 7860 2284
rect 7948 2276 7956 2284
rect 7420 2256 7428 2264
rect 7516 2256 7524 2264
rect 7580 2256 7588 2264
rect 7612 2256 7620 2264
rect 7836 2256 7844 2264
rect 7916 2256 7924 2264
rect 188 2236 196 2244
rect 204 2236 212 2244
rect 252 2236 260 2244
rect 428 2236 436 2244
rect 460 2236 468 2244
rect 620 2236 628 2244
rect 1260 2236 1268 2244
rect 1500 2236 1508 2244
rect 1852 2236 1860 2244
rect 2060 2236 2068 2244
rect 2092 2236 2100 2244
rect 2332 2236 2340 2244
rect 2572 2236 2580 2244
rect 2620 2236 2628 2244
rect 3116 2236 3124 2244
rect 3532 2236 3540 2244
rect 4124 2236 4132 2244
rect 4332 2236 4340 2244
rect 4524 2236 4532 2244
rect 4572 2236 4580 2244
rect 4892 2236 4900 2244
rect 4972 2236 4980 2244
rect 5372 2236 5380 2244
rect 5548 2236 5556 2244
rect 5692 2236 5700 2244
rect 6076 2236 6084 2244
rect 6476 2236 6484 2244
rect 6780 2236 6788 2244
rect 6828 2236 6836 2244
rect 7260 2236 7268 2244
rect 7500 2236 7508 2244
rect 7788 2236 7796 2244
rect 2316 2216 2324 2224
rect 6188 2216 6196 2224
rect 6444 2216 6452 2224
rect 7356 2216 7364 2224
rect 3278 2206 3286 2214
rect 3292 2206 3300 2214
rect 3306 2206 3314 2214
rect 6350 2206 6358 2214
rect 6364 2206 6372 2214
rect 6378 2206 6386 2214
rect 3772 2196 3780 2204
rect 4540 2196 4548 2204
rect 6988 2196 6996 2204
rect 156 2176 164 2184
rect 332 2176 340 2184
rect 524 2176 532 2184
rect 1132 2176 1140 2184
rect 1340 2176 1348 2184
rect 1372 2176 1380 2184
rect 1484 2176 1492 2184
rect 2172 2176 2180 2184
rect 2348 2176 2356 2184
rect 2540 2176 2548 2184
rect 2572 2176 2580 2184
rect 2684 2176 2692 2184
rect 2812 2176 2820 2184
rect 2860 2176 2868 2184
rect 2924 2176 2932 2184
rect 3004 2176 3012 2184
rect 3084 2176 3092 2184
rect 3148 2176 3156 2184
rect 3180 2176 3188 2184
rect 3500 2176 3508 2184
rect 3980 2176 3988 2184
rect 4012 2176 4020 2184
rect 4236 2176 4244 2184
rect 4444 2176 4452 2184
rect 4460 2176 4468 2184
rect 4524 2176 4532 2184
rect 4556 2176 4564 2184
rect 4588 2176 4596 2184
rect 4796 2176 4804 2184
rect 5340 2176 5348 2184
rect 5596 2176 5604 2184
rect 5628 2176 5636 2184
rect 5660 2176 5668 2184
rect 5884 2176 5892 2184
rect 5916 2176 5924 2184
rect 6172 2176 6180 2184
rect 6524 2176 6532 2184
rect 6604 2176 6612 2184
rect 6844 2176 6852 2184
rect 7276 2176 7284 2184
rect 7388 2176 7396 2184
rect 7580 2176 7588 2184
rect 172 2156 180 2164
rect 188 2156 196 2164
rect 716 2156 724 2164
rect 812 2156 820 2164
rect 1004 2156 1012 2164
rect 1180 2156 1188 2164
rect 1276 2156 1284 2164
rect 1500 2156 1508 2164
rect 1580 2156 1588 2164
rect 12 2136 20 2144
rect 108 2136 116 2144
rect 140 2136 148 2144
rect 284 2136 292 2144
rect 412 2136 420 2144
rect 428 2136 436 2144
rect 460 2136 468 2144
rect 476 2136 484 2144
rect 524 2136 532 2144
rect 588 2136 596 2144
rect 636 2136 644 2144
rect 732 2136 740 2144
rect 1292 2136 1300 2144
rect 1356 2136 1364 2144
rect 1388 2136 1396 2144
rect 1852 2156 1860 2164
rect 1980 2156 1988 2164
rect 2156 2156 2164 2164
rect 2700 2156 2708 2164
rect 2988 2156 2996 2164
rect 3020 2156 3028 2164
rect 3164 2156 3172 2164
rect 3692 2156 3700 2164
rect 3708 2156 3716 2164
rect 3772 2156 3780 2164
rect 3788 2156 3796 2164
rect 3900 2156 3908 2164
rect 4044 2156 4052 2164
rect 4060 2156 4068 2164
rect 4476 2156 4484 2164
rect 4540 2156 4548 2164
rect 5100 2156 5108 2164
rect 5532 2156 5540 2164
rect 5580 2156 5588 2164
rect 1708 2136 1716 2144
rect 108 2116 116 2124
rect 124 2116 132 2124
rect 236 2116 244 2124
rect 252 2116 260 2124
rect 300 2116 308 2124
rect 204 2096 212 2104
rect 268 2096 276 2104
rect 396 2116 404 2124
rect 492 2116 500 2124
rect 652 2116 660 2124
rect 668 2116 676 2124
rect 748 2116 756 2124
rect 812 2118 820 2126
rect 1020 2116 1028 2124
rect 1148 2116 1156 2124
rect 1212 2116 1220 2124
rect 1244 2116 1252 2124
rect 1308 2116 1316 2124
rect 1500 2116 1508 2124
rect 1660 2116 1668 2124
rect 1676 2116 1684 2124
rect 1788 2136 1796 2144
rect 2108 2136 2116 2144
rect 2172 2136 2180 2144
rect 2380 2136 2388 2144
rect 2572 2136 2580 2144
rect 2604 2136 2612 2144
rect 2636 2136 2644 2144
rect 2796 2136 2804 2144
rect 2844 2136 2852 2144
rect 2892 2136 2900 2144
rect 2972 2136 2980 2144
rect 3020 2136 3028 2144
rect 3132 2136 3140 2144
rect 3340 2136 3348 2144
rect 3516 2136 3524 2144
rect 3532 2136 3540 2144
rect 3628 2136 3636 2144
rect 3660 2136 3668 2144
rect 3836 2136 3844 2144
rect 3852 2136 3860 2144
rect 4028 2136 4036 2144
rect 4124 2136 4132 2144
rect 4284 2136 4292 2144
rect 4780 2136 4788 2144
rect 4988 2136 4996 2144
rect 5180 2136 5188 2144
rect 5388 2136 5396 2144
rect 5436 2136 5444 2144
rect 5468 2136 5476 2144
rect 5644 2136 5652 2144
rect 5852 2156 5860 2164
rect 6284 2156 6292 2164
rect 6364 2156 6372 2164
rect 6572 2156 6580 2164
rect 6924 2156 6932 2164
rect 6988 2156 6996 2164
rect 7292 2156 7300 2164
rect 5692 2136 5700 2144
rect 5788 2136 5796 2144
rect 5820 2136 5828 2144
rect 5868 2136 5876 2144
rect 6076 2136 6084 2144
rect 6108 2136 6116 2144
rect 6204 2136 6212 2144
rect 6220 2136 6228 2144
rect 6236 2132 6244 2140
rect 6332 2136 6340 2144
rect 6412 2136 6420 2144
rect 6444 2136 6452 2144
rect 1804 2116 1812 2124
rect 1852 2116 1860 2124
rect 1884 2116 1892 2124
rect 1932 2116 1940 2124
rect 2060 2116 2068 2124
rect 2156 2116 2164 2124
rect 2268 2116 2276 2124
rect 2316 2116 2324 2124
rect 2428 2116 2436 2124
rect 2556 2116 2564 2124
rect 2620 2116 2628 2124
rect 2652 2116 2660 2124
rect 2732 2116 2740 2124
rect 2764 2116 2772 2124
rect 2780 2116 2788 2124
rect 2924 2116 2932 2124
rect 3308 2118 3316 2126
rect 3436 2116 3444 2124
rect 3468 2116 3476 2124
rect 3596 2116 3604 2124
rect 3644 2116 3652 2124
rect 348 2096 356 2104
rect 524 2096 532 2104
rect 572 2096 580 2104
rect 668 2096 676 2104
rect 1196 2096 1204 2104
rect 1404 2096 1412 2104
rect 1436 2096 1444 2104
rect 2684 2096 2692 2104
rect 2748 2096 2756 2104
rect 2812 2096 2820 2104
rect 2860 2096 2868 2104
rect 2892 2096 2900 2104
rect 3420 2096 3428 2104
rect 3932 2116 3940 2124
rect 3948 2116 3956 2124
rect 4108 2116 4116 2124
rect 4332 2116 4340 2124
rect 4380 2116 4388 2124
rect 4492 2116 4500 2124
rect 4572 2116 4580 2124
rect 4668 2116 4676 2124
rect 4716 2118 4724 2126
rect 4956 2118 4964 2126
rect 5036 2116 5044 2124
rect 5068 2116 5076 2124
rect 5116 2116 5124 2124
rect 5260 2116 5268 2124
rect 5276 2116 5284 2124
rect 5516 2116 5524 2124
rect 5564 2116 5572 2124
rect 5724 2116 5732 2124
rect 5804 2116 5812 2124
rect 6044 2118 6052 2126
rect 6316 2116 6324 2124
rect 6460 2116 6468 2124
rect 6636 2136 6644 2144
rect 6668 2136 6676 2144
rect 6780 2136 6788 2144
rect 6796 2136 6804 2144
rect 7004 2136 7012 2144
rect 7068 2136 7076 2144
rect 7116 2136 7124 2144
rect 7148 2136 7156 2144
rect 7180 2136 7188 2144
rect 7212 2136 7220 2144
rect 7324 2136 7332 2144
rect 7372 2136 7380 2144
rect 7548 2136 7556 2144
rect 7740 2136 7748 2144
rect 7804 2136 7812 2144
rect 7820 2136 7828 2144
rect 7948 2136 7956 2144
rect 6540 2116 6548 2124
rect 6588 2116 6596 2124
rect 6652 2116 6660 2124
rect 6684 2116 6692 2124
rect 3996 2096 4004 2104
rect 5020 2096 5028 2104
rect 5356 2096 5364 2104
rect 5900 2096 5908 2104
rect 6476 2096 6484 2104
rect 6524 2096 6532 2104
rect 6716 2096 6724 2104
rect 6764 2116 6772 2124
rect 6796 2116 6804 2124
rect 6812 2116 6820 2124
rect 6892 2116 6900 2124
rect 7052 2116 7060 2124
rect 7116 2116 7124 2124
rect 7132 2116 7140 2124
rect 7212 2116 7220 2124
rect 7228 2116 7236 2124
rect 7244 2116 7252 2124
rect 7308 2116 7316 2124
rect 7500 2116 7508 2124
rect 7708 2118 7716 2126
rect 7836 2116 7844 2124
rect 7932 2118 7940 2126
rect 8076 2116 8084 2124
rect 6844 2096 6852 2104
rect 6908 2096 6916 2104
rect 7036 2096 7044 2104
rect 7260 2096 7268 2104
rect 7772 2096 7780 2104
rect 7836 2096 7844 2104
rect 7868 2096 7876 2104
rect 908 2076 916 2084
rect 940 2076 948 2084
rect 1548 2076 1556 2084
rect 1948 2076 1956 2084
rect 1980 2076 1988 2084
rect 2716 2076 2724 2084
rect 2940 2076 2948 2084
rect 3148 2076 3156 2084
rect 3372 2076 3380 2084
rect 3484 2076 3492 2084
rect 3788 2076 3796 2084
rect 3980 2076 3988 2084
rect 4060 2076 4068 2084
rect 5052 2076 5060 2084
rect 6444 2076 6452 2084
rect 6764 2076 6772 2084
rect 6876 2076 6884 2084
rect 6956 2076 6964 2084
rect 7148 2076 7156 2084
rect 7804 2076 7812 2084
rect 8060 2076 8068 2084
rect 8156 2076 8164 2084
rect 428 2036 436 2044
rect 636 2036 644 2044
rect 1596 2036 1604 2044
rect 1932 2036 1940 2044
rect 2300 2036 2308 2044
rect 3180 2036 3188 2044
rect 3692 2036 3700 2044
rect 4044 2036 4052 2044
rect 5084 2036 5092 2044
rect 5148 2036 5156 2044
rect 5500 2036 5508 2044
rect 5852 2036 5860 2044
rect 6268 2036 6276 2044
rect 6300 2036 6308 2044
rect 6892 2036 6900 2044
rect 7020 2036 7028 2044
rect 7068 2036 7076 2044
rect 7324 2036 7332 2044
rect 1742 2006 1750 2014
rect 1756 2006 1764 2014
rect 1770 2006 1778 2014
rect 4814 2006 4822 2014
rect 4828 2006 4836 2014
rect 4842 2006 4850 2014
rect 252 1976 260 1984
rect 684 1976 692 1984
rect 2620 1976 2628 1984
rect 2636 1976 2644 1984
rect 3372 1976 3380 1984
rect 3436 1976 3444 1984
rect 3500 1976 3508 1984
rect 4412 1976 4420 1984
rect 4508 1976 4516 1984
rect 4572 1976 4580 1984
rect 5052 1976 5060 1984
rect 5180 1976 5188 1984
rect 5916 1976 5924 1984
rect 6668 1976 6676 1984
rect 6748 1976 6756 1984
rect 6796 1976 6804 1984
rect 844 1956 852 1964
rect 3756 1956 3764 1964
rect 3948 1956 3956 1964
rect 7308 1956 7316 1964
rect 204 1936 212 1944
rect 668 1936 676 1944
rect 716 1936 724 1944
rect 860 1936 868 1944
rect 1020 1936 1028 1944
rect 1244 1936 1252 1944
rect 2140 1936 2148 1944
rect 2220 1936 2228 1944
rect 2972 1936 2980 1944
rect 3100 1936 3108 1944
rect 3420 1936 3428 1944
rect 3724 1936 3732 1944
rect 3820 1936 3828 1944
rect 3900 1936 3908 1944
rect 4716 1936 4724 1944
rect 5052 1936 5060 1944
rect 5324 1936 5332 1944
rect 5724 1936 5732 1944
rect 6284 1936 6292 1944
rect 7724 1936 7732 1944
rect 7948 1936 7956 1944
rect 8156 1936 8164 1944
rect 348 1916 356 1924
rect 636 1916 644 1924
rect 60 1894 68 1902
rect 204 1896 212 1904
rect 220 1896 228 1904
rect 268 1896 276 1904
rect 380 1896 388 1904
rect 492 1894 500 1902
rect 652 1896 660 1904
rect 700 1896 708 1904
rect 764 1916 772 1924
rect 828 1916 836 1924
rect 908 1916 916 1924
rect 988 1916 996 1924
rect 1212 1916 1220 1924
rect 2268 1916 2276 1924
rect 796 1896 804 1904
rect 844 1896 852 1904
rect 892 1896 900 1904
rect 1004 1896 1012 1904
rect 1068 1896 1076 1904
rect 1084 1896 1092 1904
rect 1132 1896 1140 1904
rect 1164 1896 1172 1904
rect 1196 1896 1204 1904
rect 1244 1896 1252 1904
rect 1340 1896 1348 1904
rect 1372 1896 1380 1904
rect 1404 1896 1412 1904
rect 1468 1896 1476 1904
rect 1596 1896 1604 1904
rect 1740 1896 1748 1904
rect 1788 1896 1796 1904
rect 1868 1896 1876 1904
rect 1948 1896 1956 1904
rect 1980 1896 1988 1904
rect 2124 1896 2132 1904
rect 2156 1896 2164 1904
rect 2204 1896 2212 1904
rect 2236 1896 2244 1904
rect 2396 1916 2404 1924
rect 2396 1896 2404 1904
rect 2444 1916 2452 1924
rect 2668 1916 2676 1924
rect 2748 1916 2756 1924
rect 3132 1916 3140 1924
rect 3164 1916 3172 1924
rect 3212 1916 3220 1924
rect 3228 1916 3236 1924
rect 3260 1916 3268 1924
rect 3340 1916 3348 1924
rect 3452 1916 3460 1924
rect 3836 1916 3844 1924
rect 3868 1916 3876 1924
rect 2524 1896 2532 1904
rect 2828 1896 2836 1904
rect 3020 1896 3028 1904
rect 3132 1896 3140 1904
rect 3260 1896 3268 1904
rect 3372 1896 3380 1904
rect 3436 1896 3444 1904
rect 3612 1896 3620 1904
rect 3660 1896 3668 1904
rect 3788 1896 3796 1904
rect 3836 1896 3844 1904
rect 3884 1896 3892 1904
rect 3932 1896 3940 1904
rect 3996 1916 4004 1924
rect 4092 1916 4100 1924
rect 4028 1896 4036 1904
rect 4108 1896 4116 1904
rect 4172 1896 4180 1904
rect 4188 1896 4196 1904
rect 4236 1896 4244 1904
rect 4364 1916 4372 1924
rect 4588 1916 4596 1924
rect 4956 1916 4964 1924
rect 5068 1916 5076 1924
rect 5084 1916 5092 1924
rect 5116 1916 5124 1924
rect 5148 1916 5156 1924
rect 5404 1916 5412 1924
rect 5452 1916 5460 1924
rect 5468 1916 5476 1924
rect 5660 1916 5668 1924
rect 5692 1916 5700 1924
rect 4444 1896 4452 1904
rect 4508 1896 4516 1904
rect 4620 1896 4628 1904
rect 4860 1896 4868 1904
rect 4892 1896 4900 1904
rect 4988 1896 4996 1904
rect 5052 1896 5060 1904
rect 5116 1896 5124 1904
rect 5388 1896 5396 1904
rect 5468 1896 5476 1904
rect 5500 1896 5508 1904
rect 5580 1896 5588 1904
rect 5692 1896 5700 1904
rect 5836 1896 5844 1904
rect 6028 1896 6036 1904
rect 6172 1896 6180 1904
rect 6316 1896 6324 1904
rect 6332 1896 6340 1904
rect 6412 1916 6420 1924
rect 6876 1916 6884 1924
rect 6924 1916 6932 1924
rect 7324 1916 7332 1924
rect 7500 1916 7508 1924
rect 7804 1916 7812 1924
rect 7868 1916 7876 1924
rect 6460 1896 6468 1904
rect 6492 1896 6500 1904
rect 6588 1896 6596 1904
rect 6764 1896 6772 1904
rect 6844 1896 6852 1904
rect 6988 1894 6996 1902
rect 7196 1896 7204 1904
rect 7356 1896 7364 1904
rect 7420 1896 7428 1904
rect 7452 1896 7460 1904
rect 7484 1896 7492 1904
rect 7596 1894 7604 1902
rect 7740 1896 7748 1904
rect 7772 1896 7780 1904
rect 7852 1896 7860 1904
rect 7964 1916 7972 1924
rect 8060 1916 8068 1924
rect 7916 1896 7924 1904
rect 8012 1896 8020 1904
rect 8076 1896 8084 1904
rect 92 1876 100 1884
rect 364 1876 372 1884
rect 460 1876 468 1884
rect 700 1876 708 1884
rect 812 1876 820 1884
rect 956 1876 964 1884
rect 1068 1876 1076 1884
rect 1180 1876 1188 1884
rect 1356 1876 1364 1884
rect 1420 1876 1428 1884
rect 1436 1876 1444 1884
rect 1596 1876 1604 1884
rect 1772 1876 1780 1884
rect 2188 1876 2196 1884
rect 2316 1876 2324 1884
rect 2332 1876 2340 1884
rect 2380 1876 2388 1884
rect 2492 1876 2500 1884
rect 2572 1876 2580 1884
rect 2588 1880 2596 1888
rect 2700 1876 2708 1884
rect 2748 1876 2756 1884
rect 2796 1876 2804 1884
rect 2812 1876 2820 1884
rect 2908 1876 2916 1884
rect 3004 1876 3012 1884
rect 3036 1876 3044 1884
rect 3180 1876 3188 1884
rect 3196 1876 3204 1884
rect 3276 1876 3284 1884
rect 3388 1876 3396 1884
rect 3836 1876 3844 1884
rect 3932 1876 3940 1884
rect 4060 1876 4068 1884
rect 4156 1876 4164 1884
rect 4284 1876 4292 1884
rect 4316 1876 4324 1884
rect 4396 1876 4404 1884
rect 4460 1876 4468 1884
rect 4636 1876 4644 1884
rect 4652 1876 4660 1884
rect 4764 1876 4772 1884
rect 4876 1876 4884 1884
rect 5004 1876 5012 1884
rect 5132 1876 5140 1884
rect 5196 1876 5204 1884
rect 5276 1876 5284 1884
rect 5356 1876 5364 1884
rect 5420 1876 5428 1884
rect 5564 1876 5572 1884
rect 5644 1876 5652 1884
rect 5708 1876 5716 1884
rect 5884 1876 5892 1884
rect 6012 1876 6020 1884
rect 6204 1876 6212 1884
rect 6300 1876 6308 1884
rect 6524 1876 6532 1884
rect 6556 1876 6564 1884
rect 6572 1876 6580 1884
rect 6700 1880 6708 1888
rect 6716 1876 6724 1884
rect 6860 1876 6868 1884
rect 6892 1876 6900 1884
rect 7020 1876 7028 1884
rect 7148 1876 7156 1884
rect 7340 1876 7348 1884
rect 7436 1876 7444 1884
rect 7468 1876 7476 1884
rect 7516 1876 7524 1884
rect 7532 1876 7540 1884
rect 7612 1876 7620 1884
rect 7804 1876 7812 1884
rect 7836 1876 7844 1884
rect 7852 1876 7860 1884
rect 7996 1876 8004 1884
rect 8012 1876 8020 1884
rect 8044 1876 8052 1884
rect 156 1856 164 1864
rect 268 1856 276 1864
rect 332 1856 340 1864
rect 428 1856 436 1864
rect 908 1856 916 1864
rect 940 1856 948 1864
rect 1116 1856 1124 1864
rect 1292 1856 1300 1864
rect 1676 1856 1684 1864
rect 1932 1856 1940 1864
rect 2124 1856 2132 1864
rect 2524 1856 2532 1864
rect 2556 1856 2564 1864
rect 2652 1856 2660 1864
rect 2876 1856 2884 1864
rect 3068 1856 3076 1864
rect 3084 1856 3092 1864
rect 3468 1856 3476 1864
rect 3532 1856 3540 1864
rect 3772 1856 3780 1864
rect 4220 1856 4228 1864
rect 4492 1856 4500 1864
rect 4540 1856 4548 1864
rect 4556 1856 4564 1864
rect 4764 1856 4772 1864
rect 4828 1856 4836 1864
rect 5228 1856 5236 1864
rect 5244 1856 5252 1864
rect 5340 1856 5348 1864
rect 5548 1856 5556 1864
rect 5628 1856 5636 1864
rect 6492 1856 6500 1864
rect 6588 1856 6596 1864
rect 6620 1856 6628 1864
rect 6652 1856 6660 1864
rect 6732 1856 6740 1864
rect 6780 1856 6788 1864
rect 6812 1856 6820 1864
rect 7404 1856 7412 1864
rect 620 1836 628 1844
rect 1308 1836 1316 1844
rect 1484 1836 1492 1844
rect 1692 1836 1700 1844
rect 1820 1836 1828 1844
rect 1836 1836 1844 1844
rect 2060 1836 2068 1844
rect 2076 1836 2084 1844
rect 2268 1836 2276 1844
rect 2508 1836 2516 1844
rect 2540 1836 2548 1844
rect 2732 1836 2740 1844
rect 2780 1836 2788 1844
rect 2860 1836 2868 1844
rect 2892 1836 2900 1844
rect 3052 1836 3060 1844
rect 3916 1836 3924 1844
rect 4140 1836 4148 1844
rect 4268 1836 4276 1844
rect 4412 1836 4420 1844
rect 4476 1836 4484 1844
rect 4924 1836 4932 1844
rect 5212 1836 5220 1844
rect 5260 1836 5268 1844
rect 5292 1836 5300 1844
rect 5468 1836 5476 1844
rect 5612 1836 5620 1844
rect 6476 1836 6484 1844
rect 6524 1836 6532 1844
rect 6924 1836 6932 1844
rect 7116 1836 7124 1844
rect 7820 1836 7828 1844
rect 7980 1836 7988 1844
rect 268 1816 276 1824
rect 3532 1816 3540 1824
rect 4828 1816 4836 1824
rect 3278 1806 3286 1814
rect 3292 1806 3300 1814
rect 3306 1806 3314 1814
rect 6350 1806 6358 1814
rect 6364 1806 6372 1814
rect 6378 1806 6386 1814
rect 172 1796 180 1804
rect 604 1796 612 1804
rect 5964 1796 5972 1804
rect 28 1776 36 1784
rect 588 1776 596 1784
rect 1036 1776 1044 1784
rect 1132 1776 1140 1784
rect 2188 1776 2196 1784
rect 2492 1776 2500 1784
rect 2604 1776 2612 1784
rect 2780 1776 2788 1784
rect 4060 1776 4068 1784
rect 4124 1776 4132 1784
rect 4652 1776 4660 1784
rect 4684 1776 4692 1784
rect 5084 1776 5092 1784
rect 5532 1776 5540 1784
rect 5948 1776 5956 1784
rect 6124 1776 6132 1784
rect 6140 1776 6148 1784
rect 6332 1776 6340 1784
rect 6684 1776 6692 1784
rect 6796 1776 6804 1784
rect 6844 1776 6852 1784
rect 6988 1776 6996 1784
rect 7260 1776 7268 1784
rect 7324 1776 7332 1784
rect 7564 1776 7572 1784
rect 7948 1776 7956 1784
rect 8140 1776 8148 1784
rect 156 1756 164 1764
rect 172 1756 180 1764
rect 236 1756 244 1764
rect 524 1756 532 1764
rect 540 1756 548 1764
rect 604 1756 612 1764
rect 732 1756 740 1764
rect 908 1756 916 1764
rect 924 1756 932 1764
rect 956 1756 964 1764
rect 1436 1756 1444 1764
rect 1452 1756 1460 1764
rect 1596 1756 1604 1764
rect 1660 1756 1668 1764
rect 76 1736 84 1744
rect 300 1736 308 1744
rect 636 1736 644 1744
rect 668 1736 676 1744
rect 716 1736 724 1744
rect 764 1736 772 1744
rect 796 1736 804 1744
rect 892 1736 900 1744
rect 956 1736 964 1744
rect 972 1736 980 1744
rect 1052 1736 1060 1744
rect 1068 1736 1076 1744
rect 1228 1736 1236 1744
rect 1372 1736 1380 1744
rect 1420 1736 1428 1744
rect 1836 1756 1844 1764
rect 1964 1756 1972 1764
rect 2396 1756 2404 1764
rect 2636 1756 2644 1764
rect 2684 1756 2692 1764
rect 2844 1756 2852 1764
rect 3100 1756 3108 1764
rect 3196 1756 3204 1764
rect 3212 1756 3220 1764
rect 3596 1756 3604 1764
rect 3644 1756 3652 1764
rect 3660 1756 3668 1764
rect 3804 1756 3812 1764
rect 3820 1756 3828 1764
rect 3852 1756 3860 1764
rect 4316 1756 4324 1764
rect 4700 1756 4708 1764
rect 4988 1756 4996 1764
rect 5068 1756 5076 1764
rect 5756 1756 5764 1764
rect 5964 1756 5972 1764
rect 6444 1756 6452 1764
rect 6732 1756 6740 1764
rect 6892 1756 6900 1764
rect 1868 1736 1876 1744
rect 1932 1736 1940 1744
rect 2092 1736 2100 1744
rect 2364 1736 2372 1744
rect 2428 1736 2436 1744
rect 2460 1736 2468 1744
rect 2556 1736 2564 1744
rect 2652 1736 2660 1744
rect 2700 1736 2708 1744
rect 2764 1736 2772 1744
rect 2828 1736 2836 1744
rect 2924 1736 2932 1744
rect 2940 1736 2948 1744
rect 3004 1736 3012 1744
rect 3052 1736 3060 1744
rect 3164 1736 3172 1744
rect 3276 1736 3284 1744
rect 3324 1736 3332 1744
rect 3404 1736 3412 1744
rect 3436 1736 3444 1744
rect 3500 1736 3508 1744
rect 3532 1736 3540 1744
rect 3564 1736 3572 1744
rect 3580 1736 3588 1744
rect 3724 1736 3732 1744
rect 3740 1736 3748 1744
rect 3852 1736 3860 1744
rect 3948 1736 3956 1744
rect 4012 1736 4020 1744
rect 4108 1736 4116 1744
rect 4380 1736 4388 1744
rect 4460 1736 4468 1744
rect 4492 1736 4500 1744
rect 4812 1736 4820 1744
rect 4908 1736 4916 1744
rect 5004 1736 5012 1744
rect 5084 1736 5092 1744
rect 5148 1736 5156 1744
rect 5196 1736 5204 1744
rect 5260 1736 5268 1744
rect 5292 1736 5300 1744
rect 5324 1736 5332 1744
rect 5372 1736 5380 1744
rect 5596 1736 5604 1744
rect 5628 1736 5636 1744
rect 5660 1736 5668 1744
rect 5788 1736 5796 1744
rect 6364 1736 6372 1744
rect 6508 1736 6516 1744
rect 6540 1736 6548 1744
rect 6572 1736 6580 1744
rect 6668 1736 6676 1744
rect 6748 1736 6756 1744
rect 6828 1736 6836 1744
rect 7148 1736 7156 1744
rect 7180 1736 7188 1744
rect 7276 1736 7284 1744
rect 7372 1736 7380 1744
rect 7452 1736 7460 1744
rect 7884 1736 7892 1744
rect 7980 1736 7988 1744
rect 44 1716 52 1724
rect 92 1716 100 1724
rect 108 1716 116 1724
rect 172 1716 180 1724
rect 332 1716 340 1724
rect 444 1716 452 1724
rect 476 1716 484 1724
rect 60 1696 68 1704
rect 444 1696 452 1704
rect 780 1716 788 1724
rect 796 1716 804 1724
rect 684 1696 692 1704
rect 1004 1696 1012 1704
rect 1084 1716 1092 1724
rect 1116 1716 1124 1724
rect 1260 1718 1268 1726
rect 1324 1716 1332 1724
rect 1532 1716 1540 1724
rect 1596 1718 1604 1726
rect 1692 1716 1700 1724
rect 1724 1716 1732 1724
rect 1804 1716 1812 1724
rect 1900 1718 1908 1726
rect 2092 1716 2100 1724
rect 2332 1718 2340 1726
rect 2412 1716 2420 1724
rect 2444 1716 2452 1724
rect 2588 1716 2596 1724
rect 2716 1716 2724 1724
rect 2812 1716 2820 1724
rect 2876 1716 2884 1724
rect 2956 1716 2964 1724
rect 1324 1696 1332 1704
rect 1388 1696 1396 1704
rect 1708 1696 1716 1704
rect 2076 1696 2084 1704
rect 2188 1696 2196 1704
rect 2572 1696 2580 1704
rect 2716 1696 2724 1704
rect 2748 1696 2756 1704
rect 2796 1696 2804 1704
rect 2892 1696 2900 1704
rect 3036 1716 3044 1724
rect 3068 1716 3076 1724
rect 3116 1716 3124 1724
rect 3180 1716 3188 1724
rect 3260 1716 3268 1724
rect 3356 1716 3364 1724
rect 3212 1696 3220 1704
rect 3404 1716 3412 1724
rect 3436 1716 3444 1724
rect 3500 1716 3508 1724
rect 3516 1716 3524 1724
rect 3580 1716 3588 1724
rect 3628 1716 3636 1724
rect 3676 1716 3684 1724
rect 3756 1716 3764 1724
rect 3404 1696 3412 1704
rect 3756 1696 3764 1704
rect 3788 1696 3796 1704
rect 3820 1696 3828 1704
rect 3900 1696 3908 1704
rect 3996 1716 4004 1724
rect 4028 1716 4036 1724
rect 4076 1716 4084 1724
rect 4188 1716 4196 1724
rect 4252 1718 4260 1726
rect 4364 1716 4372 1724
rect 4444 1716 4452 1724
rect 4524 1718 4532 1726
rect 4668 1716 4676 1724
rect 4828 1716 4836 1724
rect 5244 1716 5252 1724
rect 5276 1716 5284 1724
rect 5340 1716 5348 1724
rect 5404 1718 5412 1726
rect 4396 1696 4404 1704
rect 4412 1696 4420 1704
rect 5212 1696 5220 1704
rect 5228 1696 5236 1704
rect 5628 1716 5636 1724
rect 5708 1716 5716 1724
rect 5724 1716 5732 1724
rect 5820 1718 5828 1726
rect 6076 1716 6084 1724
rect 6204 1716 6212 1724
rect 6236 1716 6244 1724
rect 6460 1716 6468 1724
rect 6492 1716 6500 1724
rect 6524 1716 6532 1724
rect 6588 1716 6596 1724
rect 6620 1716 6628 1724
rect 5596 1696 5604 1704
rect 6332 1696 6340 1704
rect 6604 1696 6612 1704
rect 6780 1696 6788 1704
rect 6876 1716 6884 1724
rect 6924 1716 6932 1724
rect 6972 1716 6980 1724
rect 7084 1716 7092 1724
rect 7228 1716 7236 1724
rect 6972 1696 6980 1704
rect 7308 1696 7316 1704
rect 7356 1716 7364 1724
rect 7436 1718 7444 1726
rect 7644 1716 7652 1724
rect 7708 1718 7716 1726
rect 7820 1718 7828 1726
rect 8012 1718 8020 1726
rect 28 1676 36 1684
rect 156 1676 164 1684
rect 1164 1676 1172 1684
rect 2156 1676 2164 1684
rect 2204 1676 2212 1684
rect 2604 1676 2612 1684
rect 2668 1676 2676 1684
rect 2988 1676 2996 1684
rect 3452 1676 3460 1684
rect 4444 1676 4452 1684
rect 4748 1676 4756 1684
rect 4988 1676 4996 1684
rect 5036 1676 5044 1684
rect 6636 1676 6644 1684
rect 6700 1676 6708 1684
rect 7212 1676 7220 1684
rect 7612 1676 7620 1684
rect 7580 1656 7588 1664
rect 428 1636 436 1644
rect 732 1636 740 1644
rect 1468 1636 1476 1644
rect 1676 1636 1684 1644
rect 3132 1636 3140 1644
rect 3356 1636 3364 1644
rect 3532 1636 3540 1644
rect 3724 1636 3732 1644
rect 3932 1636 3940 1644
rect 3964 1636 3972 1644
rect 4716 1636 4724 1644
rect 5292 1636 5300 1644
rect 5692 1636 5700 1644
rect 5980 1636 5988 1644
rect 6044 1636 6052 1644
rect 6380 1636 6388 1644
rect 6572 1636 6580 1644
rect 6620 1636 6628 1644
rect 7196 1636 7204 1644
rect 7260 1636 7268 1644
rect 1742 1606 1750 1614
rect 1756 1606 1764 1614
rect 1770 1606 1778 1614
rect 4814 1606 4822 1614
rect 4828 1606 4836 1614
rect 4842 1606 4850 1614
rect 44 1576 52 1584
rect 92 1576 100 1584
rect 940 1576 948 1584
rect 1452 1576 1460 1584
rect 1644 1576 1652 1584
rect 2348 1576 2356 1584
rect 2540 1576 2548 1584
rect 2780 1576 2788 1584
rect 2796 1576 2804 1584
rect 3020 1576 3028 1584
rect 3212 1576 3220 1584
rect 4076 1576 4084 1584
rect 4652 1576 4660 1584
rect 4780 1576 4788 1584
rect 5932 1576 5940 1584
rect 6236 1576 6244 1584
rect 7100 1576 7108 1584
rect 7404 1576 7412 1584
rect 7708 1576 7716 1584
rect 1948 1556 1956 1564
rect 4044 1556 4052 1564
rect 5276 1556 5284 1564
rect 5708 1556 5716 1564
rect 6940 1556 6948 1564
rect 28 1536 36 1544
rect 44 1536 52 1544
rect 460 1536 468 1544
rect 1132 1536 1140 1544
rect 1228 1536 1236 1544
rect 1340 1536 1348 1544
rect 1548 1536 1556 1544
rect 3596 1536 3604 1544
rect 3740 1536 3748 1544
rect 4012 1536 4020 1544
rect 4204 1536 4212 1544
rect 4252 1536 4260 1544
rect 5724 1536 5732 1544
rect 6124 1536 6132 1544
rect 6252 1536 6260 1544
rect 6860 1536 6868 1544
rect 7724 1536 7732 1544
rect 7772 1536 7780 1544
rect 7900 1536 7908 1544
rect 76 1516 84 1524
rect 108 1516 116 1524
rect 172 1516 180 1524
rect 236 1516 244 1524
rect 44 1496 52 1504
rect 124 1496 132 1504
rect 140 1496 148 1504
rect 316 1496 324 1504
rect 396 1496 404 1504
rect 428 1496 436 1504
rect 444 1496 452 1504
rect 1164 1516 1172 1524
rect 1196 1516 1204 1524
rect 1580 1516 1588 1524
rect 1628 1516 1636 1524
rect 1756 1516 1764 1524
rect 1836 1516 1844 1524
rect 2252 1516 2260 1524
rect 3228 1516 3236 1524
rect 4140 1516 4148 1524
rect 540 1496 548 1504
rect 572 1496 580 1504
rect 620 1496 628 1504
rect 764 1494 772 1502
rect 828 1496 836 1504
rect 908 1496 916 1504
rect 1020 1496 1028 1504
rect 1068 1496 1076 1504
rect 1148 1496 1156 1504
rect 1228 1496 1236 1504
rect 1356 1496 1364 1504
rect 1404 1496 1412 1504
rect 1468 1496 1476 1504
rect 1516 1496 1524 1504
rect 1564 1496 1572 1504
rect 1692 1496 1700 1504
rect 1708 1496 1716 1504
rect 1772 1496 1780 1504
rect 1884 1496 1892 1504
rect 2076 1496 2084 1504
rect 2172 1496 2180 1504
rect 2284 1496 2292 1504
rect 2300 1496 2308 1504
rect 2316 1496 2324 1504
rect 2412 1494 2420 1502
rect 2668 1496 2676 1504
rect 2716 1496 2724 1504
rect 2828 1496 2836 1504
rect 2908 1496 2916 1504
rect 3100 1496 3108 1504
rect 3260 1496 3268 1504
rect 3420 1494 3428 1502
rect 3676 1496 3684 1504
rect 3932 1496 3940 1504
rect 4204 1496 4212 1504
rect 4316 1516 4324 1524
rect 4364 1516 4372 1524
rect 5228 1516 5236 1524
rect 5260 1516 5268 1524
rect 5548 1516 5556 1524
rect 5612 1516 5620 1524
rect 5692 1516 5700 1524
rect 5820 1516 5828 1524
rect 5852 1516 5860 1524
rect 6156 1516 6164 1524
rect 6284 1516 6292 1524
rect 6396 1516 6404 1524
rect 6540 1516 6548 1524
rect 6780 1516 6788 1524
rect 7084 1516 7092 1524
rect 7628 1516 7636 1524
rect 7692 1516 7700 1524
rect 7804 1516 7812 1524
rect 7820 1516 7828 1524
rect 7932 1516 7940 1524
rect 7964 1516 7972 1524
rect 4284 1496 4292 1504
rect 4348 1496 4356 1504
rect 4396 1496 4404 1504
rect 4524 1494 4532 1502
rect 4588 1496 4596 1504
rect 4700 1496 4708 1504
rect 4732 1496 4740 1504
rect 4812 1496 4820 1504
rect 4892 1496 4900 1504
rect 4940 1496 4948 1504
rect 5116 1494 5124 1502
rect 5228 1496 5236 1504
rect 5340 1496 5348 1504
rect 5404 1494 5412 1502
rect 5484 1496 5492 1504
rect 5708 1496 5716 1504
rect 5756 1496 5764 1504
rect 5820 1496 5828 1504
rect 5868 1496 5876 1504
rect 5884 1496 5892 1504
rect 6092 1496 6100 1504
rect 6108 1496 6116 1504
rect 6172 1496 6180 1504
rect 6268 1496 6276 1504
rect 6300 1496 6308 1504
rect 6508 1496 6516 1504
rect 6620 1496 6628 1504
rect 6652 1496 6660 1504
rect 6876 1496 6884 1504
rect 6908 1496 6916 1504
rect 6988 1496 6996 1504
rect 7052 1496 7060 1504
rect 7084 1496 7092 1504
rect 7180 1496 7188 1504
rect 7196 1496 7204 1504
rect 7436 1496 7444 1504
rect 7500 1496 7508 1504
rect 7708 1496 7716 1504
rect 7772 1496 7780 1504
rect 7852 1496 7860 1504
rect 7900 1496 7908 1504
rect 156 1476 164 1484
rect 220 1476 228 1484
rect 268 1476 276 1484
rect 332 1476 340 1484
rect 348 1476 356 1484
rect 412 1476 420 1484
rect 492 1476 500 1484
rect 524 1476 532 1484
rect 540 1476 548 1484
rect 636 1476 644 1484
rect 684 1480 692 1488
rect 700 1476 708 1484
rect 972 1476 980 1484
rect 1148 1476 1156 1484
rect 1212 1476 1220 1484
rect 1292 1476 1300 1484
rect 1340 1476 1348 1484
rect 1404 1476 1412 1484
rect 1596 1476 1604 1484
rect 1676 1476 1684 1484
rect 1692 1476 1700 1484
rect 1868 1476 1876 1484
rect 1916 1476 1924 1484
rect 2012 1476 2020 1484
rect 2060 1476 2068 1484
rect 2172 1476 2180 1484
rect 2220 1476 2228 1484
rect 2380 1476 2388 1484
rect 2556 1476 2564 1484
rect 2588 1476 2596 1484
rect 2620 1476 2628 1484
rect 2860 1476 2868 1484
rect 3052 1476 3060 1484
rect 3244 1476 3252 1484
rect 3388 1476 3396 1484
rect 3564 1476 3572 1484
rect 3628 1476 3636 1484
rect 3692 1476 3700 1484
rect 3772 1476 3780 1484
rect 3884 1476 3892 1484
rect 4060 1476 4068 1484
rect 4108 1476 4116 1484
rect 4172 1476 4180 1484
rect 4188 1476 4196 1484
rect 4300 1476 4308 1484
rect 4316 1476 4324 1484
rect 4364 1476 4372 1484
rect 4396 1476 4404 1484
rect 4716 1476 4724 1484
rect 4876 1476 4884 1484
rect 5052 1476 5060 1484
rect 5100 1476 5108 1484
rect 5436 1476 5444 1484
rect 5468 1476 5476 1484
rect 5580 1476 5588 1484
rect 5628 1476 5636 1484
rect 5660 1476 5668 1484
rect 5836 1476 5844 1484
rect 5900 1476 5908 1484
rect 6108 1476 6116 1484
rect 6188 1476 6196 1484
rect 6380 1476 6388 1484
rect 6444 1476 6452 1484
rect 6540 1476 6548 1484
rect 6780 1476 6788 1484
rect 6812 1476 6820 1484
rect 6860 1476 6868 1484
rect 6988 1476 6996 1484
rect 7292 1476 7300 1484
rect 7468 1476 7476 1484
rect 7484 1476 7492 1484
rect 7756 1476 7764 1484
rect 7868 1476 7876 1484
rect 7884 1476 7892 1484
rect 8012 1476 8020 1484
rect 8156 1476 8164 1484
rect 76 1456 84 1464
rect 284 1456 292 1464
rect 572 1456 580 1464
rect 1228 1456 1236 1464
rect 1308 1456 1316 1464
rect 1484 1456 1492 1464
rect 1644 1456 1652 1464
rect 1900 1456 1908 1464
rect 2044 1456 2052 1464
rect 2268 1456 2276 1464
rect 3356 1456 3364 1464
rect 3788 1456 3796 1464
rect 3852 1456 3860 1464
rect 4428 1456 4436 1464
rect 4444 1456 4452 1464
rect 4620 1456 4628 1464
rect 4764 1456 4772 1464
rect 4972 1456 4980 1464
rect 5180 1456 5188 1464
rect 5340 1456 5348 1464
rect 5564 1456 5572 1464
rect 5772 1456 5780 1464
rect 6220 1456 6228 1464
rect 6460 1456 6468 1464
rect 6748 1456 6756 1464
rect 6908 1456 6916 1464
rect 7004 1456 7012 1464
rect 7548 1456 7556 1464
rect 7580 1456 7588 1464
rect 7644 1456 7652 1464
rect 7660 1456 7668 1464
rect 7964 1456 7972 1464
rect 7996 1456 8004 1464
rect 172 1436 180 1444
rect 348 1436 356 1444
rect 492 1436 500 1444
rect 652 1436 660 1444
rect 892 1436 900 1444
rect 1388 1436 1396 1444
rect 1564 1436 1572 1444
rect 1628 1436 1636 1444
rect 2028 1436 2036 1444
rect 2108 1436 2116 1444
rect 2124 1436 2132 1444
rect 2188 1436 2196 1444
rect 2796 1436 2804 1444
rect 3548 1436 3556 1444
rect 3692 1436 3700 1444
rect 3804 1436 3812 1444
rect 4460 1436 4468 1444
rect 4668 1436 4676 1444
rect 4748 1436 4756 1444
rect 4780 1436 4788 1444
rect 4924 1436 4932 1444
rect 4956 1436 4964 1444
rect 4988 1436 4996 1444
rect 6060 1436 6068 1444
rect 6204 1436 6212 1444
rect 6556 1436 6564 1444
rect 7532 1436 7540 1444
rect 7564 1436 7572 1444
rect 7676 1436 7684 1444
rect 7820 1436 7828 1444
rect 7948 1436 7956 1444
rect 8044 1436 8052 1444
rect 3788 1416 3796 1424
rect 7644 1416 7652 1424
rect 3278 1406 3286 1414
rect 3292 1406 3300 1414
rect 3306 1406 3314 1414
rect 6350 1406 6358 1414
rect 6364 1406 6372 1414
rect 6378 1406 6386 1414
rect 668 1396 676 1404
rect 5948 1396 5956 1404
rect 380 1376 388 1384
rect 428 1376 436 1384
rect 524 1376 532 1384
rect 556 1376 564 1384
rect 1052 1376 1060 1384
rect 1100 1376 1108 1384
rect 1180 1376 1188 1384
rect 1260 1376 1268 1384
rect 1308 1376 1316 1384
rect 1532 1376 1540 1384
rect 2140 1376 2148 1384
rect 2492 1376 2500 1384
rect 2908 1376 2916 1384
rect 3724 1376 3732 1384
rect 3836 1376 3844 1384
rect 3916 1376 3924 1384
rect 3980 1376 3988 1384
rect 4044 1376 4052 1384
rect 4092 1376 4100 1384
rect 4428 1376 4436 1384
rect 5388 1376 5396 1384
rect 5564 1376 5572 1384
rect 5596 1376 5604 1384
rect 5692 1376 5700 1384
rect 5852 1376 5860 1384
rect 5932 1376 5940 1384
rect 5964 1376 5972 1384
rect 6124 1376 6132 1384
rect 6668 1376 6676 1384
rect 7116 1376 7124 1384
rect 7756 1376 7764 1384
rect 7836 1376 7844 1384
rect 172 1356 180 1364
rect 444 1356 452 1364
rect 604 1356 612 1364
rect 668 1356 676 1364
rect 1084 1356 1092 1364
rect 1164 1356 1172 1364
rect 1340 1356 1348 1364
rect 1852 1356 1860 1364
rect 2060 1356 2068 1364
rect 2252 1356 2260 1364
rect 2300 1356 2308 1364
rect 2332 1356 2340 1364
rect 2620 1356 2628 1364
rect 2876 1356 2884 1364
rect 3532 1356 3540 1364
rect 3596 1356 3604 1364
rect 3820 1356 3828 1364
rect 3900 1356 3908 1364
rect 3932 1356 3940 1364
rect 12 1336 20 1344
rect 108 1336 116 1344
rect 140 1336 148 1344
rect 412 1336 420 1344
rect 460 1336 468 1344
rect 556 1336 564 1344
rect 588 1336 596 1344
rect 1004 1336 1012 1344
rect 1020 1336 1028 1344
rect 1148 1336 1156 1344
rect 1196 1336 1204 1344
rect 1276 1336 1284 1344
rect 1324 1336 1332 1344
rect 1420 1336 1428 1344
rect 1484 1336 1492 1344
rect 1500 1336 1508 1344
rect 1612 1336 1620 1344
rect 1644 1336 1652 1344
rect 1916 1336 1924 1344
rect 1964 1336 1972 1344
rect 1980 1336 1988 1344
rect 2028 1336 2036 1344
rect 2108 1336 2116 1344
rect 2156 1336 2164 1344
rect 2188 1336 2196 1344
rect 2364 1336 2372 1344
rect 2460 1336 2468 1344
rect 2860 1336 2868 1344
rect 2892 1336 2900 1344
rect 3068 1336 3076 1344
rect 3100 1336 3108 1344
rect 3212 1336 3220 1344
rect 3452 1336 3460 1344
rect 3500 1336 3508 1344
rect 3516 1336 3524 1344
rect 3740 1336 3748 1344
rect 3884 1336 3892 1344
rect 4764 1356 4772 1364
rect 4780 1356 4788 1364
rect 4908 1356 4916 1364
rect 4956 1356 4964 1364
rect 5196 1356 5204 1364
rect 5276 1356 5284 1364
rect 5308 1356 5316 1364
rect 5484 1356 5492 1364
rect 5548 1356 5556 1364
rect 5612 1356 5620 1364
rect 5628 1356 5636 1364
rect 5724 1356 5732 1364
rect 5740 1356 5748 1364
rect 5868 1356 5876 1364
rect 5884 1356 5892 1364
rect 5948 1356 5956 1364
rect 7308 1356 7316 1364
rect 7708 1356 7716 1364
rect 7900 1356 7908 1364
rect 4012 1336 4020 1344
rect 4076 1336 4084 1344
rect 4108 1336 4116 1344
rect 4268 1336 4276 1344
rect 4332 1336 4340 1344
rect 4396 1336 4404 1344
rect 4508 1336 4516 1344
rect 4620 1336 4628 1344
rect 4716 1336 4724 1344
rect 4876 1336 4884 1344
rect 5052 1336 5060 1344
rect 5276 1336 5284 1344
rect 5324 1336 5332 1344
rect 5436 1336 5444 1344
rect 5452 1336 5460 1344
rect 5500 1336 5508 1344
rect 5772 1336 5780 1344
rect 5788 1332 5796 1340
rect 6156 1336 6164 1344
rect 6236 1336 6244 1344
rect 6460 1336 6468 1344
rect 6572 1336 6580 1344
rect 6588 1336 6596 1344
rect 6684 1336 6692 1344
rect 6796 1336 6804 1344
rect 6908 1336 6916 1344
rect 6972 1336 6980 1344
rect 7356 1336 7364 1344
rect 7452 1336 7460 1344
rect 7532 1336 7540 1344
rect 7580 1336 7588 1344
rect 7596 1336 7604 1344
rect 7628 1336 7636 1344
rect 7692 1336 7700 1344
rect 7804 1336 7812 1344
rect 7852 1336 7860 1344
rect 7948 1336 7956 1344
rect 7980 1336 7988 1344
rect 44 1316 52 1324
rect 124 1316 132 1324
rect 172 1316 180 1324
rect 236 1318 244 1326
rect 300 1316 308 1324
rect 380 1296 388 1304
rect 492 1296 500 1304
rect 668 1316 676 1324
rect 748 1316 756 1324
rect 796 1316 804 1324
rect 876 1316 884 1324
rect 1132 1316 1140 1324
rect 556 1296 564 1304
rect 1052 1296 1060 1304
rect 1228 1296 1236 1304
rect 1372 1316 1380 1324
rect 1436 1316 1444 1324
rect 1468 1316 1476 1324
rect 1580 1316 1588 1324
rect 1628 1316 1636 1324
rect 1852 1318 1860 1326
rect 1948 1316 1956 1324
rect 2076 1316 2084 1324
rect 2172 1316 2180 1324
rect 2236 1316 2244 1324
rect 2332 1316 2340 1324
rect 2412 1316 2420 1324
rect 2620 1318 2628 1326
rect 2684 1316 2692 1324
rect 3036 1318 3044 1326
rect 3116 1316 3124 1324
rect 3132 1316 3140 1324
rect 3228 1316 3236 1324
rect 3356 1316 3364 1324
rect 3628 1316 3636 1324
rect 3788 1316 3796 1324
rect 3868 1316 3876 1324
rect 3964 1316 3972 1324
rect 4060 1316 4068 1324
rect 4124 1316 4132 1324
rect 4172 1316 4180 1324
rect 4220 1316 4228 1324
rect 4284 1316 4292 1324
rect 4348 1316 4356 1324
rect 4380 1316 4388 1324
rect 4604 1316 4612 1324
rect 4716 1316 4724 1324
rect 4732 1316 4740 1324
rect 4860 1316 4868 1324
rect 4908 1316 4916 1324
rect 4924 1316 4932 1324
rect 5020 1318 5028 1326
rect 5164 1316 5172 1324
rect 5196 1316 5204 1324
rect 5244 1316 5252 1324
rect 5276 1316 5284 1324
rect 5436 1316 5444 1324
rect 5468 1316 5476 1324
rect 5580 1316 5588 1324
rect 5692 1316 5700 1324
rect 5756 1316 5764 1324
rect 5996 1316 6004 1324
rect 6220 1318 6228 1326
rect 6412 1316 6420 1324
rect 6476 1316 6484 1324
rect 1404 1296 1412 1304
rect 1436 1296 1444 1304
rect 1596 1296 1604 1304
rect 1660 1296 1668 1304
rect 1916 1296 1924 1304
rect 2060 1296 2068 1304
rect 2396 1296 2404 1304
rect 3148 1296 3156 1304
rect 3404 1296 3412 1304
rect 3468 1296 3476 1304
rect 3740 1296 3748 1304
rect 4044 1296 4052 1304
rect 4188 1296 4196 1304
rect 4204 1296 4212 1304
rect 4316 1296 4324 1304
rect 4348 1296 4356 1304
rect 4380 1296 4388 1304
rect 4460 1296 4468 1304
rect 4524 1296 4532 1304
rect 5532 1296 5540 1304
rect 5644 1296 5652 1304
rect 5708 1296 5716 1304
rect 6508 1296 6516 1304
rect 6556 1316 6564 1324
rect 6636 1316 6644 1324
rect 6700 1316 6708 1324
rect 6780 1316 6788 1324
rect 6924 1316 6932 1324
rect 7100 1316 7108 1324
rect 7180 1316 7188 1324
rect 7244 1318 7252 1326
rect 7404 1316 7412 1324
rect 7756 1316 7764 1324
rect 7916 1316 7924 1324
rect 7948 1316 7956 1324
rect 8012 1318 8020 1326
rect 6620 1296 6628 1304
rect 7532 1296 7540 1304
rect 7628 1296 7636 1304
rect 7740 1296 7748 1304
rect 7836 1296 7844 1304
rect 7884 1296 7892 1304
rect 364 1276 372 1284
rect 1276 1276 1284 1284
rect 1468 1276 1476 1284
rect 1532 1276 1540 1284
rect 1564 1276 1572 1284
rect 1724 1276 1732 1284
rect 1980 1276 1988 1284
rect 2124 1276 2132 1284
rect 4156 1276 4164 1284
rect 4220 1276 4228 1284
rect 4236 1276 4244 1284
rect 4556 1276 4564 1284
rect 5676 1276 5684 1284
rect 6892 1276 6900 1284
rect 6956 1276 6964 1284
rect 7516 1276 7524 1284
rect 7644 1276 7652 1284
rect 7772 1276 7780 1284
rect 4284 1256 4292 1264
rect 860 1236 868 1244
rect 1068 1236 1076 1244
rect 1580 1236 1588 1244
rect 2044 1236 2052 1244
rect 2220 1236 2228 1244
rect 2348 1236 2356 1244
rect 2428 1236 2436 1244
rect 2716 1236 2724 1244
rect 2844 1236 2852 1244
rect 3388 1236 3396 1244
rect 4252 1236 4260 1244
rect 4748 1236 4756 1244
rect 4940 1236 4948 1244
rect 5148 1236 5156 1244
rect 5164 1236 5172 1244
rect 5516 1236 5524 1244
rect 6348 1236 6356 1244
rect 6444 1236 6452 1244
rect 6556 1236 6564 1244
rect 6924 1236 6932 1244
rect 7324 1236 7332 1244
rect 7868 1236 7876 1244
rect 8140 1236 8148 1244
rect 1742 1206 1750 1214
rect 1756 1206 1764 1214
rect 1770 1206 1778 1214
rect 4814 1206 4822 1214
rect 4828 1206 4836 1214
rect 4842 1206 4850 1214
rect 364 1176 372 1184
rect 748 1176 756 1184
rect 1820 1176 1828 1184
rect 2044 1176 2052 1184
rect 2668 1176 2676 1184
rect 3196 1176 3204 1184
rect 3276 1176 3284 1184
rect 3436 1176 3444 1184
rect 3564 1176 3572 1184
rect 3756 1176 3764 1184
rect 3980 1176 3988 1184
rect 4236 1176 4244 1184
rect 4492 1176 4500 1184
rect 5068 1176 5076 1184
rect 5212 1176 5220 1184
rect 6892 1176 6900 1184
rect 7084 1176 7092 1184
rect 7100 1176 7108 1184
rect 7244 1176 7252 1184
rect 7340 1176 7348 1184
rect 3068 1156 3076 1164
rect 5340 1156 5348 1164
rect 764 1136 772 1144
rect 860 1136 868 1144
rect 2476 1136 2484 1144
rect 2620 1136 2628 1144
rect 2684 1136 2692 1144
rect 3404 1136 3412 1144
rect 3772 1136 3780 1144
rect 4524 1136 4532 1144
rect 5052 1136 5060 1144
rect 5404 1136 5412 1144
rect 6604 1136 6612 1144
rect 6620 1136 6628 1144
rect 6748 1136 6756 1144
rect 6844 1136 6852 1144
rect 6860 1136 6868 1144
rect 7516 1136 7524 1144
rect 8156 1136 8164 1144
rect 460 1116 468 1124
rect 668 1116 676 1124
rect 732 1116 740 1124
rect 124 1096 132 1104
rect 348 1096 356 1104
rect 396 1096 404 1104
rect 428 1096 436 1104
rect 556 1096 564 1104
rect 572 1096 580 1104
rect 700 1096 708 1104
rect 748 1096 756 1104
rect 860 1096 868 1104
rect 908 1116 916 1124
rect 988 1116 996 1124
rect 940 1096 948 1104
rect 1116 1096 1124 1104
rect 1244 1116 1252 1124
rect 1436 1116 1444 1124
rect 1548 1116 1556 1124
rect 1708 1116 1716 1124
rect 1324 1096 1332 1104
rect 1356 1096 1364 1104
rect 2316 1116 2324 1124
rect 2396 1116 2404 1124
rect 2412 1116 2420 1124
rect 2508 1116 2516 1124
rect 2572 1116 2580 1124
rect 1932 1096 1940 1104
rect 2092 1096 2100 1104
rect 2140 1096 2148 1104
rect 2204 1096 2212 1104
rect 2364 1096 2372 1104
rect 2412 1096 2420 1104
rect 2492 1096 2500 1104
rect 172 1076 180 1084
rect 204 1076 212 1084
rect 300 1076 308 1084
rect 412 1076 420 1084
rect 716 1076 724 1084
rect 796 1076 804 1084
rect 844 1076 852 1084
rect 956 1076 964 1084
rect 1036 1076 1044 1084
rect 1164 1076 1172 1084
rect 1196 1076 1204 1084
rect 1276 1076 1284 1084
rect 1340 1076 1348 1084
rect 1404 1076 1412 1084
rect 1564 1076 1572 1084
rect 1660 1076 1668 1084
rect 1676 1076 1684 1084
rect 1756 1076 1764 1084
rect 1804 1076 1812 1084
rect 1980 1076 1988 1084
rect 2140 1076 2148 1084
rect 2156 1076 2164 1084
rect 2204 1076 2212 1084
rect 2300 1076 2308 1084
rect 2348 1076 2356 1084
rect 2380 1076 2388 1084
rect 2444 1076 2452 1084
rect 2540 1096 2548 1104
rect 2652 1116 2660 1124
rect 2796 1116 2804 1124
rect 3388 1116 3396 1124
rect 3628 1116 3636 1124
rect 4044 1116 4052 1124
rect 4732 1116 4740 1124
rect 4764 1116 4772 1124
rect 4908 1116 4916 1124
rect 4956 1116 4964 1124
rect 4988 1116 4996 1124
rect 5084 1116 5092 1124
rect 5244 1116 5252 1124
rect 5260 1116 5268 1124
rect 5292 1116 5300 1124
rect 5372 1116 5380 1124
rect 5708 1116 5716 1124
rect 5724 1116 5732 1124
rect 5772 1116 5780 1124
rect 5868 1116 5876 1124
rect 5900 1116 5908 1124
rect 5916 1116 5924 1124
rect 6076 1116 6084 1124
rect 6236 1116 6244 1124
rect 6268 1116 6276 1124
rect 6700 1116 6708 1124
rect 6748 1116 6756 1124
rect 6796 1116 6804 1124
rect 6812 1116 6820 1124
rect 7180 1116 7188 1124
rect 7196 1116 7204 1124
rect 7212 1116 7220 1124
rect 7308 1116 7316 1124
rect 7372 1116 7380 1124
rect 7612 1116 7620 1124
rect 2620 1096 2628 1104
rect 2668 1096 2676 1104
rect 2732 1096 2740 1104
rect 2812 1096 2820 1104
rect 2828 1096 2836 1104
rect 2940 1094 2948 1102
rect 3228 1096 3236 1104
rect 3292 1096 3300 1104
rect 3436 1096 3444 1104
rect 3500 1096 3508 1104
rect 3548 1096 3556 1104
rect 3660 1096 3668 1104
rect 3884 1096 3892 1104
rect 3964 1096 3972 1104
rect 4028 1096 4036 1104
rect 4140 1096 4148 1104
rect 4284 1096 4292 1104
rect 4348 1094 4356 1102
rect 4588 1096 4596 1104
rect 4652 1094 4660 1102
rect 4732 1096 4740 1104
rect 4764 1096 4772 1104
rect 5004 1096 5012 1104
rect 5068 1096 5076 1104
rect 5116 1096 5124 1104
rect 5212 1096 5220 1104
rect 5244 1096 5252 1104
rect 5340 1096 5348 1104
rect 5388 1096 5396 1104
rect 5532 1096 5540 1104
rect 5676 1096 5684 1104
rect 5708 1096 5716 1104
rect 5788 1096 5796 1104
rect 5932 1096 5940 1104
rect 5980 1096 5988 1104
rect 6028 1096 6036 1104
rect 6092 1096 6100 1104
rect 6156 1096 6164 1104
rect 6188 1096 6196 1104
rect 6220 1096 6228 1104
rect 6268 1096 6276 1104
rect 6364 1096 6372 1104
rect 6476 1094 6484 1102
rect 6652 1096 6660 1104
rect 6764 1096 6772 1104
rect 6828 1096 6836 1104
rect 6956 1094 6964 1102
rect 7132 1096 7140 1104
rect 7244 1096 7252 1104
rect 2636 1076 2644 1084
rect 2908 1076 2916 1084
rect 3084 1076 3092 1084
rect 3228 1076 3236 1084
rect 3276 1076 3284 1084
rect 3356 1076 3364 1084
rect 3372 1076 3380 1084
rect 3452 1076 3460 1084
rect 3596 1076 3604 1084
rect 3660 1076 3668 1084
rect 3708 1076 3716 1084
rect 3724 1080 3732 1088
rect 3932 1076 3940 1084
rect 3980 1076 3988 1084
rect 4012 1076 4020 1084
rect 4076 1080 4084 1088
rect 4092 1076 4100 1084
rect 988 1056 996 1064
rect 1020 1056 1028 1064
rect 1036 1056 1044 1064
rect 1100 1056 1108 1064
rect 1452 1056 1460 1064
rect 1500 1056 1508 1064
rect 2012 1056 2020 1064
rect 2076 1056 2084 1064
rect 2188 1056 2196 1064
rect 2332 1056 2340 1064
rect 2492 1056 2500 1064
rect 2716 1056 2724 1064
rect 2780 1056 2788 1064
rect 2876 1056 2884 1064
rect 3468 1056 3476 1064
rect 3532 1056 3540 1064
rect 3692 1056 3700 1064
rect 4140 1076 4148 1084
rect 4236 1076 4244 1084
rect 4268 1076 4276 1084
rect 4716 1076 4724 1084
rect 4892 1080 4900 1088
rect 7420 1096 7428 1104
rect 7484 1096 7492 1104
rect 8140 1116 8148 1124
rect 7660 1096 7668 1104
rect 7852 1096 7860 1104
rect 7932 1096 7940 1104
rect 7980 1096 7988 1104
rect 4908 1076 4916 1084
rect 4988 1076 4996 1084
rect 5020 1076 5028 1084
rect 5100 1076 5108 1084
rect 5148 1076 5156 1084
rect 5292 1076 5300 1084
rect 5356 1076 5364 1084
rect 5420 1076 5428 1084
rect 5756 1076 5764 1084
rect 5820 1076 5828 1084
rect 5916 1076 5924 1084
rect 5948 1076 5956 1084
rect 6044 1076 6052 1084
rect 6172 1076 6180 1084
rect 6204 1076 6212 1084
rect 6444 1076 6452 1084
rect 6620 1076 6628 1084
rect 6668 1076 6676 1084
rect 6732 1076 6740 1084
rect 6924 1076 6932 1084
rect 7148 1076 7156 1084
rect 7356 1076 7364 1084
rect 7372 1076 7380 1084
rect 7420 1076 7428 1084
rect 7436 1076 7444 1084
rect 7452 1076 7460 1084
rect 7468 1076 7476 1084
rect 7532 1076 7540 1084
rect 7564 1076 7572 1084
rect 7676 1076 7684 1084
rect 7756 1076 7764 1084
rect 7868 1076 7876 1084
rect 7900 1076 7908 1084
rect 8028 1076 8036 1084
rect 8060 1076 8068 1084
rect 8108 1076 8116 1084
rect 4140 1056 4148 1064
rect 4204 1056 4212 1064
rect 4348 1056 4356 1064
rect 4508 1056 4516 1064
rect 4796 1056 4804 1064
rect 5180 1056 5188 1064
rect 5564 1056 5572 1064
rect 5628 1056 5636 1064
rect 5852 1056 5860 1064
rect 6108 1056 6116 1064
rect 6316 1056 6324 1064
rect 6332 1056 6340 1064
rect 6876 1056 6884 1064
rect 7276 1056 7284 1064
rect 7500 1056 7508 1064
rect 7548 1056 7556 1064
rect 7708 1056 7716 1064
rect 7772 1056 7780 1064
rect 7820 1056 7828 1064
rect 7964 1056 7972 1064
rect 12 1036 20 1044
rect 236 1036 244 1044
rect 316 1036 324 1044
rect 460 1036 468 1044
rect 652 1036 660 1044
rect 668 1036 676 1044
rect 812 1036 820 1044
rect 972 1036 980 1044
rect 1132 1036 1140 1044
rect 1292 1036 1300 1044
rect 1388 1036 1396 1044
rect 1420 1036 1428 1044
rect 1468 1036 1476 1044
rect 1484 1036 1492 1044
rect 1532 1036 1540 1044
rect 1596 1036 1604 1044
rect 1740 1036 1748 1044
rect 2172 1036 2180 1044
rect 4188 1036 4196 1044
rect 4476 1036 4484 1044
rect 4812 1036 4820 1044
rect 5436 1036 5444 1044
rect 5708 1036 5716 1044
rect 6012 1036 6020 1044
rect 6348 1036 6356 1044
rect 6700 1036 6708 1044
rect 7372 1036 7380 1044
rect 7628 1036 7636 1044
rect 7724 1036 7732 1044
rect 7788 1036 7796 1044
rect 7884 1036 7892 1044
rect 7996 1036 8004 1044
rect 2076 1016 2084 1024
rect 2716 1016 2724 1024
rect 7772 1016 7780 1024
rect 3278 1006 3286 1014
rect 3292 1006 3300 1014
rect 3306 1006 3314 1014
rect 6350 1006 6358 1014
rect 6364 1006 6372 1014
rect 6378 1006 6386 1014
rect 2460 996 2468 1004
rect 5148 996 5156 1004
rect 6460 996 6468 1004
rect 124 976 132 984
rect 572 976 580 984
rect 780 976 788 984
rect 1820 976 1828 984
rect 2012 976 2020 984
rect 2252 976 2260 984
rect 2908 976 2916 984
rect 3516 976 3524 984
rect 3564 976 3572 984
rect 3628 976 3636 984
rect 3740 976 3748 984
rect 3836 976 3844 984
rect 4220 976 4228 984
rect 4380 976 4388 984
rect 4460 976 4468 984
rect 4732 976 4740 984
rect 4876 976 4884 984
rect 5004 976 5012 984
rect 5068 976 5076 984
rect 5164 976 5172 984
rect 5228 976 5236 984
rect 5596 976 5604 984
rect 5628 976 5636 984
rect 6892 976 6900 984
rect 6908 976 6916 984
rect 7036 976 7044 984
rect 7468 976 7476 984
rect 7900 976 7908 984
rect 8140 976 8148 984
rect 12 956 20 964
rect 140 956 148 964
rect 236 956 244 964
rect 508 956 516 964
rect 540 956 548 964
rect 556 956 564 964
rect 636 956 644 964
rect 1212 956 1220 964
rect 1548 956 1556 964
rect 1804 956 1812 964
rect 2460 956 2468 964
rect 2524 956 2532 964
rect 2700 956 2708 964
rect 2716 956 2724 964
rect 2924 956 2932 964
rect 3180 956 3188 964
rect 3212 956 3220 964
rect 3228 956 3236 964
rect 3692 956 3700 964
rect 3852 956 3860 964
rect 4204 956 4212 964
rect 4508 956 4516 964
rect 4988 956 4996 964
rect 5020 956 5028 964
rect 5052 956 5060 964
rect 5148 956 5156 964
rect 5212 956 5220 964
rect 5740 956 5748 964
rect 6268 956 6276 964
rect 6396 956 6404 964
rect 6460 956 6468 964
rect 6924 956 6932 964
rect 7740 956 7748 964
rect 7804 956 7812 964
rect 44 936 52 944
rect 108 936 116 944
rect 156 936 164 944
rect 188 936 196 944
rect 300 936 308 944
rect 364 936 372 944
rect 588 936 596 944
rect 652 936 660 944
rect 748 936 756 944
rect 828 936 836 944
rect 956 936 964 944
rect 1068 936 1076 944
rect 1116 936 1124 944
rect 1180 936 1188 944
rect 1276 936 1284 944
rect 1292 936 1300 944
rect 1340 936 1348 944
rect 1404 936 1412 944
rect 1484 936 1492 944
rect 1580 936 1588 944
rect 1612 936 1620 944
rect 1708 936 1716 944
rect 1980 936 1988 944
rect 2124 936 2132 944
rect 2204 936 2212 944
rect 2428 936 2436 944
rect 2540 936 2548 944
rect 2620 936 2628 944
rect 2636 936 2644 944
rect 2716 936 2724 944
rect 2956 936 2964 944
rect 3068 936 3076 944
rect 3132 936 3140 944
rect 3196 936 3204 944
rect 3228 936 3236 944
rect 3260 936 3268 944
rect 3404 936 3412 944
rect 3612 936 3620 944
rect 3708 936 3716 944
rect 3788 936 3796 944
rect 3804 936 3812 944
rect 3948 936 3956 944
rect 4060 936 4068 944
rect 4268 936 4276 944
rect 4316 936 4324 944
rect 4412 936 4420 944
rect 4428 936 4436 944
rect 4588 936 4596 944
rect 4604 936 4612 944
rect 4684 936 4692 944
rect 4860 936 4868 944
rect 4892 936 4900 944
rect 4924 936 4932 944
rect 5084 936 5092 944
rect 5388 936 5396 944
rect 5612 936 5620 944
rect 5772 936 5780 944
rect 6124 936 6132 944
rect 6204 936 6212 944
rect 6380 936 6388 944
rect 6476 936 6484 944
rect 6572 936 6580 944
rect 6604 936 6612 944
rect 6700 936 6708 944
rect 6780 936 6788 944
rect 6940 936 6948 944
rect 7004 936 7012 944
rect 7276 936 7284 944
rect 7356 936 7364 944
rect 7404 936 7412 944
rect 7436 936 7444 944
rect 7596 936 7604 944
rect 7644 936 7652 944
rect 8012 936 8020 944
rect 8092 936 8100 944
rect 92 916 100 924
rect 172 916 180 924
rect 204 916 212 924
rect 300 916 308 924
rect 364 916 372 924
rect 412 916 420 924
rect 444 916 452 924
rect 780 916 788 924
rect 876 916 884 924
rect 908 916 916 924
rect 940 916 948 924
rect 972 916 980 924
rect 60 896 68 904
rect 76 896 84 904
rect 204 896 212 904
rect 316 896 324 904
rect 428 896 436 904
rect 764 896 772 904
rect 860 896 868 904
rect 1036 916 1044 924
rect 1116 916 1124 924
rect 1164 916 1172 924
rect 1260 916 1268 924
rect 1308 916 1316 924
rect 1372 916 1380 924
rect 1388 916 1396 924
rect 1436 916 1444 924
rect 1500 916 1508 924
rect 1564 916 1572 924
rect 1596 916 1604 924
rect 1660 916 1668 924
rect 1724 916 1732 924
rect 1932 916 1940 924
rect 2140 918 2148 926
rect 2220 916 2228 924
rect 2396 918 2404 926
rect 1084 896 1092 904
rect 1132 896 1140 904
rect 1228 896 1236 904
rect 1260 896 1268 904
rect 1340 896 1348 904
rect 1356 896 1364 904
rect 1420 896 1428 904
rect 1644 896 1652 904
rect 2572 896 2580 904
rect 2636 916 2644 924
rect 2684 916 2692 924
rect 2780 918 2788 926
rect 2844 916 2852 924
rect 2972 916 2980 924
rect 2684 896 2692 904
rect 3004 896 3012 904
rect 3052 916 3060 924
rect 3292 916 3300 924
rect 3356 916 3364 924
rect 3548 916 3556 924
rect 3596 916 3604 924
rect 3660 916 3668 924
rect 3116 896 3124 904
rect 3180 896 3188 904
rect 3340 896 3348 904
rect 3644 896 3652 904
rect 3916 916 3924 924
rect 3964 916 3972 924
rect 3756 896 3764 904
rect 3836 896 3844 904
rect 3932 896 3940 904
rect 3996 896 4004 904
rect 4044 916 4052 924
rect 4108 916 4116 924
rect 4140 916 4148 924
rect 4268 916 4276 924
rect 4476 916 4484 924
rect 4524 916 4532 924
rect 4556 916 4564 924
rect 4124 896 4132 904
rect 4300 896 4308 904
rect 4460 896 4468 904
rect 4700 916 4708 924
rect 4780 916 4788 924
rect 4908 916 4916 924
rect 4972 916 4980 924
rect 5100 916 5108 924
rect 5356 918 5364 926
rect 5484 916 5492 924
rect 5532 916 5540 924
rect 5676 916 5684 924
rect 5708 916 5716 924
rect 5804 918 5812 926
rect 5868 916 5876 924
rect 5980 916 5988 924
rect 5996 916 6004 924
rect 6172 916 6180 924
rect 6300 916 6308 924
rect 6588 916 6596 924
rect 6652 916 6660 924
rect 6684 916 6692 924
rect 6764 918 6772 926
rect 7052 916 7060 924
rect 7068 916 7076 924
rect 7244 918 7252 926
rect 7340 916 7348 924
rect 7404 916 7412 924
rect 8108 932 8116 940
rect 7516 916 7524 924
rect 7564 916 7572 924
rect 7580 916 7588 924
rect 7740 918 7748 926
rect 7852 916 7860 924
rect 8028 918 8036 926
rect 4652 896 4660 904
rect 4748 896 4756 904
rect 4924 896 4932 904
rect 5644 896 5652 904
rect 5660 896 5668 904
rect 6172 896 6180 904
rect 6236 896 6244 904
rect 6284 896 6292 904
rect 6444 896 6452 904
rect 6652 896 6660 904
rect 6972 896 6980 904
rect 7308 896 7316 904
rect 7404 896 7412 904
rect 7468 896 7476 904
rect 7548 896 7556 904
rect 7852 896 7860 904
rect 7884 896 7892 904
rect 284 876 292 884
rect 348 876 356 884
rect 396 876 404 884
rect 636 876 644 884
rect 684 876 692 884
rect 796 876 804 884
rect 1004 876 1012 884
rect 1452 876 1460 884
rect 1532 876 1540 884
rect 1756 876 1764 884
rect 3292 876 3300 884
rect 3372 876 3380 884
rect 3436 876 3444 884
rect 3900 876 3908 884
rect 4044 876 4052 884
rect 4092 876 4100 884
rect 4844 876 4852 884
rect 5020 876 5028 884
rect 5932 876 5940 884
rect 6140 876 6148 884
rect 6540 876 6548 884
rect 7388 876 7396 884
rect 7500 876 7508 884
rect 3868 856 3876 864
rect 3916 856 3924 864
rect 7484 856 7492 864
rect 28 836 36 844
rect 412 836 420 844
rect 524 836 532 844
rect 1436 836 1444 844
rect 1500 836 1508 844
rect 1676 836 1684 844
rect 2268 836 2276 844
rect 2476 836 2484 844
rect 2604 836 2612 844
rect 3052 836 3060 844
rect 3356 836 3364 844
rect 4108 836 4116 844
rect 4284 836 4292 844
rect 4780 836 4788 844
rect 5132 836 5140 844
rect 5948 836 5956 844
rect 7116 836 7124 844
rect 7340 836 7348 844
rect 7612 836 7620 844
rect 7900 836 7908 844
rect 8140 836 8148 844
rect 1742 806 1750 814
rect 1756 806 1764 814
rect 1770 806 1778 814
rect 4814 806 4822 814
rect 4828 806 4836 814
rect 4842 806 4850 814
rect 268 776 276 784
rect 588 776 596 784
rect 604 776 612 784
rect 1004 776 1012 784
rect 1212 776 1220 784
rect 1340 776 1348 784
rect 2044 776 2052 784
rect 2172 776 2180 784
rect 2396 776 2404 784
rect 2636 776 2644 784
rect 2748 776 2756 784
rect 3836 776 3844 784
rect 4108 776 4116 784
rect 4540 776 4548 784
rect 4556 776 4564 784
rect 4988 776 4996 784
rect 5868 776 5876 784
rect 7020 776 7028 784
rect 7468 776 7476 784
rect 7756 776 7764 784
rect 8044 776 8052 784
rect 284 736 292 744
rect 1228 736 1236 744
rect 1372 736 1380 744
rect 2380 736 2388 744
rect 2940 736 2948 744
rect 3340 736 3348 744
rect 5132 736 5140 744
rect 5228 736 5236 744
rect 5564 736 5572 744
rect 7004 736 7012 744
rect 7180 736 7188 744
rect 8060 736 8068 744
rect 60 716 68 724
rect 28 696 36 704
rect 140 716 148 724
rect 252 716 260 724
rect 316 716 324 724
rect 1372 716 1380 724
rect 1580 716 1588 724
rect 1772 716 1780 724
rect 2220 716 2228 724
rect 2284 716 2292 724
rect 172 696 180 704
rect 300 696 308 704
rect 332 696 340 704
rect 396 696 404 704
rect 460 694 468 702
rect 684 694 692 702
rect 908 696 916 704
rect 1116 696 1124 704
rect 1388 696 1396 704
rect 1548 696 1556 704
rect 1628 696 1636 704
rect 1644 696 1652 704
rect 1676 696 1684 704
rect 1708 696 1716 704
rect 1788 696 1796 704
rect 1804 696 1812 704
rect 1916 694 1924 702
rect 1980 696 1988 704
rect 2252 696 2260 704
rect 2332 716 2340 724
rect 2412 716 2420 724
rect 2476 716 2484 724
rect 2828 716 2836 724
rect 2924 716 2932 724
rect 3372 716 3380 724
rect 3612 716 3620 724
rect 3708 716 3716 724
rect 3852 716 3860 724
rect 4140 716 4148 724
rect 4156 716 4164 724
rect 4268 716 4276 724
rect 5068 716 5076 724
rect 5100 716 5108 724
rect 2332 696 2340 704
rect 2396 696 2404 704
rect 2444 696 2452 704
rect 2476 696 2484 704
rect 2588 696 2596 704
rect 2604 696 2612 704
rect 2684 696 2692 704
rect 2700 696 2708 704
rect 2764 696 2772 704
rect 2796 696 2804 704
rect 2844 696 2852 704
rect 2876 696 2884 704
rect 3004 696 3012 704
rect 3036 696 3044 704
rect 3356 696 3364 704
rect 3388 696 3396 704
rect 3516 694 3524 702
rect 3692 696 3700 704
rect 3788 696 3796 704
rect 3884 696 3892 704
rect 4012 696 4020 704
rect 4108 696 4116 704
rect 4140 696 4148 704
rect 4236 696 4244 704
rect 4284 696 4292 704
rect 4316 696 4324 704
rect 4412 694 4420 702
rect 4684 694 4692 702
rect 4844 694 4852 702
rect 5036 696 5044 704
rect 5100 696 5108 704
rect 5516 716 5524 724
rect 5532 716 5540 724
rect 5180 696 5188 704
rect 5212 696 5220 704
rect 5340 696 5348 704
rect 5420 696 5428 704
rect 12 676 20 684
rect 92 676 100 684
rect 124 676 132 684
rect 172 676 180 684
rect 220 676 228 684
rect 252 676 260 684
rect 348 676 356 684
rect 380 676 388 684
rect 396 676 404 684
rect 492 676 500 684
rect 700 676 708 684
rect 844 676 852 684
rect 1036 676 1044 684
rect 1116 676 1124 684
rect 1292 676 1300 684
rect 1436 676 1444 684
rect 1452 680 1460 688
rect 1692 676 1700 684
rect 1884 676 1892 684
rect 2060 676 2068 684
rect 2236 676 2244 684
rect 2348 676 2356 684
rect 2428 676 2436 684
rect 2492 676 2500 684
rect 2556 676 2564 684
rect 2620 676 2628 684
rect 2668 676 2676 684
rect 2716 676 2724 684
rect 2748 676 2756 684
rect 2780 676 2788 684
rect 2924 676 2932 684
rect 3132 676 3140 684
rect 3260 676 3268 684
rect 3340 676 3348 684
rect 3484 676 3492 684
rect 3740 676 3748 684
rect 3804 676 3812 684
rect 3900 676 3908 684
rect 3932 676 3940 684
rect 3980 676 3988 684
rect 4076 676 4084 684
rect 4092 676 4100 684
rect 4188 676 4196 684
rect 4300 676 4308 684
rect 4380 676 4388 684
rect 4876 676 4884 684
rect 5020 676 5028 684
rect 5068 676 5076 684
rect 5084 676 5092 684
rect 5148 676 5156 684
rect 5196 676 5204 684
rect 5388 676 5396 684
rect 5436 680 5444 688
rect 5564 696 5572 704
rect 5644 694 5652 702
rect 5692 696 5700 704
rect 5804 696 5812 704
rect 5852 696 5860 704
rect 5980 716 5988 724
rect 6428 716 6436 724
rect 6476 716 6484 724
rect 6012 696 6020 704
rect 6540 716 6548 724
rect 7356 716 7364 724
rect 7372 716 7380 724
rect 7596 716 7604 724
rect 7852 716 7860 724
rect 7980 716 7988 724
rect 8028 716 8036 724
rect 8108 716 8116 724
rect 8156 716 8164 724
rect 6140 694 6148 702
rect 6652 696 6660 704
rect 6812 696 6820 704
rect 6876 694 6884 702
rect 7052 696 7060 704
rect 7116 696 7124 704
rect 7164 696 7172 704
rect 7244 696 7252 704
rect 7324 696 7332 704
rect 7420 696 7428 704
rect 7788 696 7796 704
rect 8044 696 8052 704
rect 8108 696 8116 704
rect 5484 676 5492 684
rect 5580 676 5588 684
rect 5788 676 5796 684
rect 5868 676 5876 684
rect 5900 676 5908 684
rect 5932 676 5940 684
rect 6012 676 6020 684
rect 6156 676 6164 684
rect 6316 680 6324 688
rect 6332 676 6340 684
rect 6444 676 6452 684
rect 6492 676 6500 684
rect 620 656 628 664
rect 1228 656 1236 664
rect 1292 656 1300 664
rect 1500 656 1508 664
rect 1596 656 1604 664
rect 1852 656 1860 664
rect 1980 656 1988 664
rect 6620 676 6628 684
rect 6716 676 6724 684
rect 6732 676 6740 684
rect 6780 676 6788 684
rect 6844 676 6852 684
rect 7068 676 7076 684
rect 7212 676 7220 684
rect 7372 676 7380 684
rect 7404 676 7412 684
rect 7452 676 7460 684
rect 7516 676 7524 684
rect 7548 676 7556 684
rect 7676 676 7684 684
rect 7836 676 7844 684
rect 7868 676 7876 684
rect 7964 676 7972 684
rect 8012 676 8020 684
rect 8092 676 8100 684
rect 2204 656 2212 664
rect 2556 656 2564 664
rect 2572 656 2580 664
rect 2844 656 2852 664
rect 3452 656 3460 664
rect 3516 656 3524 664
rect 3820 656 3828 664
rect 3964 656 3972 664
rect 4252 656 4260 664
rect 4684 656 4692 664
rect 5004 656 5012 664
rect 6060 656 6068 664
rect 6412 656 6420 664
rect 6588 656 6596 664
rect 6748 656 6756 664
rect 6812 656 6820 664
rect 7260 656 7268 664
rect 7276 656 7284 664
rect 7484 656 7492 664
rect 7548 656 7556 664
rect 7676 656 7684 664
rect 7724 656 7732 664
rect 7740 656 7748 664
rect 7772 656 7780 664
rect 7836 656 7844 664
rect 348 636 356 644
rect 812 636 820 644
rect 1196 636 1204 644
rect 1244 636 1252 644
rect 1388 636 1396 644
rect 1484 636 1492 644
rect 1580 636 1588 644
rect 2476 636 2484 644
rect 3644 636 3652 644
rect 3660 636 3668 644
rect 3708 636 3716 644
rect 3756 636 3764 644
rect 3852 636 3860 644
rect 3948 636 3956 644
rect 4348 636 4356 644
rect 4972 636 4980 644
rect 5516 636 5524 644
rect 5772 636 5780 644
rect 5836 636 5844 644
rect 6076 636 6084 644
rect 6268 636 6276 644
rect 6284 636 6292 644
rect 6460 636 6468 644
rect 6508 636 6516 644
rect 6604 636 6612 644
rect 7084 636 7092 644
rect 7132 636 7140 644
rect 7356 636 7364 644
rect 7532 636 7540 644
rect 7932 636 7940 644
rect 7980 636 7988 644
rect 7740 616 7748 624
rect 3278 606 3286 614
rect 3292 606 3300 614
rect 3306 606 3314 614
rect 6350 606 6358 614
rect 6364 606 6372 614
rect 6378 606 6386 614
rect 1324 596 1332 604
rect 2764 596 2772 604
rect 3196 596 3204 604
rect 6876 596 6884 604
rect 7196 596 7204 604
rect 12 576 20 584
rect 300 576 308 584
rect 1036 576 1044 584
rect 1244 576 1252 584
rect 1516 576 1524 584
rect 1676 576 1684 584
rect 2188 576 2196 584
rect 2252 576 2260 584
rect 2316 576 2324 584
rect 2380 576 2388 584
rect 2636 576 2644 584
rect 2668 576 2676 584
rect 2860 576 2868 584
rect 2892 576 2900 584
rect 3436 576 3444 584
rect 3628 576 3636 584
rect 3740 576 3748 584
rect 3932 576 3940 584
rect 4252 576 4260 584
rect 4780 576 4788 584
rect 4908 576 4916 584
rect 5036 576 5044 584
rect 5132 576 5140 584
rect 5228 576 5236 584
rect 5452 576 5460 584
rect 5708 576 5716 584
rect 5804 576 5812 584
rect 6860 576 6868 584
rect 7276 576 7284 584
rect 7468 576 7476 584
rect 7516 576 7524 584
rect 8092 576 8100 584
rect 332 556 340 564
rect 364 556 372 564
rect 476 556 484 564
rect 572 556 580 564
rect 1116 556 1124 564
rect 1260 556 1268 564
rect 1324 556 1332 564
rect 1564 556 1572 564
rect 1868 556 1876 564
rect 1932 556 1940 564
rect 2060 556 2068 564
rect 2236 556 2244 564
rect 2444 556 2452 564
rect 2716 556 2724 564
rect 2748 556 2756 564
rect 2764 556 2772 564
rect 2812 556 2820 564
rect 3132 556 3140 564
rect 3196 556 3204 564
rect 3644 556 3652 564
rect 4124 556 4132 564
rect 4268 556 4276 564
rect 4892 556 4900 564
rect 4924 556 4932 564
rect 4956 556 4964 564
rect 4988 556 4996 564
rect 5468 556 5476 564
rect 5772 556 5780 564
rect 5820 556 5828 564
rect 5852 556 5860 564
rect 6188 556 6196 564
rect 6300 556 6308 564
rect 6316 556 6324 564
rect 6540 556 6548 564
rect 6556 556 6564 564
rect 6876 556 6884 564
rect 6940 556 6948 564
rect 7196 556 7204 564
rect 7260 556 7268 564
rect 172 536 180 544
rect 204 536 212 544
rect 252 536 260 544
rect 284 536 292 544
rect 428 536 436 544
rect 924 536 932 544
rect 1388 536 1396 544
rect 1532 536 1540 544
rect 1580 536 1588 544
rect 1644 536 1652 544
rect 1900 536 1908 544
rect 1996 536 2004 544
rect 2108 536 2116 544
rect 2124 536 2132 544
rect 8060 556 8068 564
rect 2268 536 2276 544
rect 2284 532 2292 540
rect 2412 536 2420 544
rect 2476 536 2484 544
rect 2652 536 2660 544
rect 2844 536 2852 544
rect 3068 536 3076 544
rect 3340 536 3348 544
rect 3516 536 3524 544
rect 4028 536 4036 544
rect 4220 536 4228 544
rect 4284 536 4292 544
rect 4300 536 4308 544
rect 4348 536 4356 544
rect 4396 536 4404 544
rect 4684 536 4692 544
rect 5004 536 5012 544
rect 5052 536 5060 544
rect 5148 536 5156 544
rect 5180 536 5188 544
rect 5260 536 5268 544
rect 5612 536 5620 544
rect 5628 536 5636 544
rect 5724 536 5732 544
rect 6060 536 6068 544
rect 6092 536 6100 544
rect 6220 536 6228 544
rect 6236 536 6244 544
rect 6268 536 6276 544
rect 6412 536 6420 544
rect 6460 536 6468 544
rect 6572 536 6580 544
rect 6684 536 6692 544
rect 6764 536 6772 544
rect 6812 536 6820 544
rect 7020 536 7028 544
rect 7116 536 7124 544
rect 7132 536 7140 544
rect 7436 536 7444 544
rect 7500 536 7508 544
rect 7932 536 7940 544
rect 8060 536 8068 544
rect 8140 536 8148 544
rect 92 516 100 524
rect 380 516 388 524
rect 412 516 420 524
rect 444 516 452 524
rect 524 516 532 524
rect 636 518 644 526
rect 700 516 708 524
rect 780 516 788 524
rect 1148 516 1156 524
rect 1404 516 1412 524
rect 1644 516 1652 524
rect 1868 518 1876 526
rect 1980 516 1988 524
rect 2028 516 2036 524
rect 2076 516 2084 524
rect 2348 516 2356 524
rect 2396 516 2404 524
rect 2508 518 2516 526
rect 2572 516 2580 524
rect 2732 516 2740 524
rect 2924 516 2932 524
rect 3084 516 3092 524
rect 3340 516 3348 524
rect 3516 516 3524 524
rect 3692 516 3700 524
rect 3708 516 3716 524
rect 3804 516 3812 524
rect 3868 518 3876 526
rect 4060 518 4068 526
rect 4172 516 4180 524
rect 4188 516 4196 524
rect 4508 516 4516 524
rect 4668 516 4676 524
rect 4796 516 4804 524
rect 4988 516 4996 524
rect 5100 516 5108 524
rect 252 496 260 504
rect 492 496 500 504
rect 524 496 532 504
rect 1564 496 1572 504
rect 1676 496 1684 504
rect 2012 496 2020 504
rect 2332 496 2340 504
rect 2444 496 2452 504
rect 2684 496 2692 504
rect 2876 496 2884 504
rect 3724 496 3732 504
rect 4204 496 4212 504
rect 4268 496 4276 504
rect 4332 496 4340 504
rect 4396 496 4404 504
rect 5036 496 5044 504
rect 5084 496 5092 504
rect 5212 496 5220 504
rect 5340 516 5348 524
rect 5388 516 5396 524
rect 5516 516 5524 524
rect 5532 516 5540 524
rect 5596 516 5604 524
rect 5676 516 5684 524
rect 5740 516 5748 524
rect 5788 516 5796 524
rect 5932 516 5940 524
rect 5964 516 5972 524
rect 6076 516 6084 524
rect 5564 496 5572 504
rect 5660 496 5668 504
rect 6156 516 6164 524
rect 6220 516 6228 524
rect 6252 516 6260 524
rect 6284 516 6292 524
rect 6332 516 6340 524
rect 6396 516 6404 524
rect 6460 516 6468 524
rect 6508 516 6516 524
rect 6524 496 6532 504
rect 6620 496 6628 504
rect 6668 516 6676 524
rect 6732 516 6740 524
rect 6860 516 6868 524
rect 6988 516 6996 524
rect 7036 516 7044 524
rect 7052 516 7060 524
rect 6748 496 6756 504
rect 6796 496 6804 504
rect 7340 516 7348 524
rect 7356 516 7364 524
rect 7580 516 7588 524
rect 7628 516 7636 524
rect 7772 516 7780 524
rect 7964 516 7972 524
rect 8028 516 8036 524
rect 8124 516 8132 524
rect 7004 496 7012 504
rect 7068 496 7076 504
rect 7084 496 7092 504
rect 7180 496 7188 504
rect 7996 496 8004 504
rect 8092 496 8100 504
rect 1644 476 1652 484
rect 1692 476 1700 484
rect 2364 476 2372 484
rect 2812 476 2820 484
rect 6044 476 6052 484
rect 6124 476 6132 484
rect 6492 476 6500 484
rect 6668 476 6676 484
rect 6716 476 6724 484
rect 6988 476 6996 484
rect 7468 476 7476 484
rect 8060 476 8068 484
rect 6508 456 6516 464
rect 460 436 468 444
rect 764 436 772 444
rect 1036 436 1044 444
rect 1308 436 1316 444
rect 2060 436 2068 444
rect 2700 436 2708 444
rect 2956 436 2964 444
rect 3116 436 3124 444
rect 3180 436 3188 444
rect 3436 436 3444 444
rect 4412 436 4420 444
rect 4940 436 4948 444
rect 5836 436 5844 444
rect 6444 436 6452 444
rect 6700 436 6708 444
rect 6956 436 6964 444
rect 7148 436 7156 444
rect 7884 436 7892 444
rect 7916 436 7924 444
rect 1742 406 1750 414
rect 1756 406 1764 414
rect 1770 406 1778 414
rect 4814 406 4822 414
rect 4828 406 4836 414
rect 4842 406 4850 414
rect 1132 376 1140 384
rect 1228 376 1236 384
rect 1836 376 1844 384
rect 2908 376 2916 384
rect 3260 376 3268 384
rect 3340 376 3348 384
rect 4348 376 4356 384
rect 4508 376 4516 384
rect 4700 376 4708 384
rect 5100 376 5108 384
rect 5420 376 5428 384
rect 5644 376 5652 384
rect 5692 376 5700 384
rect 6396 376 6404 384
rect 6972 376 6980 384
rect 7452 376 7460 384
rect 7580 376 7588 384
rect 348 356 356 364
rect 1564 356 1572 364
rect 3020 356 3028 364
rect 3676 356 3684 364
rect 3804 356 3812 364
rect 4636 356 4644 364
rect 5228 356 5236 364
rect 220 336 228 344
rect 364 336 372 344
rect 620 336 628 344
rect 1580 336 1588 344
rect 1740 336 1748 344
rect 2444 336 2452 344
rect 2860 336 2868 344
rect 2924 336 2932 344
rect 3356 336 3364 344
rect 3548 336 3556 344
rect 3692 336 3700 344
rect 3964 336 3972 344
rect 4236 336 4244 344
rect 4428 336 4436 344
rect 4620 336 4628 344
rect 4684 336 4692 344
rect 5068 336 5076 344
rect 5116 336 5124 344
rect 5244 336 5252 344
rect 5580 336 5588 344
rect 5980 356 5988 364
rect 7020 356 7028 364
rect 5644 336 5652 344
rect 5660 336 5668 344
rect 5740 336 5748 344
rect 6956 336 6964 344
rect 252 316 260 324
rect 316 316 324 324
rect 332 316 340 324
rect 444 316 452 324
rect 492 316 500 324
rect 508 316 516 324
rect 588 316 596 324
rect 860 316 868 324
rect 1548 316 1556 324
rect 1676 316 1684 324
rect 1708 316 1716 324
rect 1932 316 1940 324
rect 2412 316 2420 324
rect 2476 316 2484 324
rect 2588 316 2596 324
rect 2604 316 2612 324
rect 2700 316 2708 324
rect 140 294 148 302
rect 204 296 212 304
rect 236 296 244 304
rect 284 296 292 304
rect 348 296 356 304
rect 396 296 404 304
rect 460 296 468 304
rect 540 296 548 304
rect 572 296 580 304
rect 716 294 724 302
rect 780 296 788 304
rect 876 296 884 304
rect 892 296 900 304
rect 1004 294 1012 302
rect 1244 296 1252 304
rect 1420 296 1428 304
rect 1564 296 1572 304
rect 1676 296 1684 304
rect 1740 296 1748 304
rect 1820 296 1828 304
rect 2012 296 2020 304
rect 2076 294 2084 302
rect 2204 296 2212 304
rect 2380 296 2388 304
rect 2396 296 2404 304
rect 2524 296 2532 304
rect 2556 296 2564 304
rect 2668 296 2676 304
rect 2748 316 2756 324
rect 2780 316 2788 324
rect 2812 316 2820 324
rect 2892 316 2900 324
rect 3292 316 3300 324
rect 3388 316 3396 324
rect 3484 316 3492 324
rect 2748 296 2756 304
rect 2844 296 2852 304
rect 2908 296 2916 304
rect 2956 296 2964 304
rect 3004 296 3012 304
rect 3068 296 3076 304
rect 3132 294 3140 302
rect 3340 296 3348 304
rect 3420 296 3428 304
rect 3484 296 3492 304
rect 3548 296 3556 304
rect 3596 316 3604 324
rect 3660 316 3668 324
rect 3900 316 3908 324
rect 3932 316 3940 324
rect 3628 296 3636 304
rect 3676 296 3684 304
rect 3724 296 3732 304
rect 3772 296 3780 304
rect 3868 296 3876 304
rect 3916 296 3924 304
rect 4588 316 4596 324
rect 4652 316 4660 324
rect 4716 316 4724 324
rect 5020 316 5028 324
rect 4044 296 4052 304
rect 4108 294 4116 302
rect 4252 296 4260 304
rect 4300 296 4308 304
rect 4364 296 4372 304
rect 4428 296 4436 304
rect 4444 296 4452 304
rect 4460 296 4468 304
rect 4476 296 4484 304
rect 4556 296 4564 304
rect 4636 296 4644 304
rect 4700 296 4708 304
rect 4988 296 4996 304
rect 5148 316 5156 324
rect 5164 316 5172 324
rect 5196 316 5204 324
rect 5612 316 5620 324
rect 5628 316 5636 324
rect 5772 316 5780 324
rect 5804 316 5812 324
rect 5836 316 5844 324
rect 5852 316 5860 324
rect 5916 316 5924 324
rect 6252 316 6260 324
rect 6892 316 6900 324
rect 6988 316 6996 324
rect 7084 316 7092 324
rect 7692 316 7700 324
rect 7708 316 7716 324
rect 7756 316 7764 324
rect 7852 316 7860 324
rect 7868 316 7876 324
rect 5068 296 5076 304
rect 5132 296 5140 304
rect 5228 296 5236 304
rect 5276 296 5284 304
rect 172 276 180 284
rect 268 276 276 284
rect 476 276 484 284
rect 556 276 564 284
rect 620 276 628 284
rect 1036 276 1044 284
rect 1148 276 1156 284
rect 1244 276 1252 284
rect 1340 276 1348 284
rect 1372 276 1380 284
rect 1692 276 1700 284
rect 1756 276 1764 284
rect 1804 276 1812 284
rect 1868 276 1876 284
rect 1884 276 1892 284
rect 2156 276 2164 284
rect 2476 276 2484 284
rect 2508 276 2516 284
rect 2540 276 2548 284
rect 2572 276 2580 284
rect 2636 276 2644 284
rect 2764 276 2772 284
rect 2812 276 2820 284
rect 2876 276 2884 284
rect 3052 276 3060 284
rect 3100 276 3108 284
rect 3164 276 3172 284
rect 3484 276 3492 284
rect 3532 276 3540 284
rect 3644 276 3652 284
rect 316 256 324 264
rect 396 256 404 264
rect 428 256 436 264
rect 524 256 532 264
rect 652 256 660 264
rect 940 256 948 264
rect 1068 256 1076 264
rect 1196 256 1204 264
rect 1612 256 1620 264
rect 1628 256 1636 264
rect 3756 276 3764 284
rect 3900 276 3908 284
rect 3916 276 3924 284
rect 3980 276 3988 284
rect 4028 276 4036 284
rect 4124 276 4132 284
rect 4172 276 4180 284
rect 4316 276 4324 284
rect 4492 276 4500 284
rect 4508 276 4516 284
rect 4540 276 4548 284
rect 4732 276 4740 284
rect 4828 276 4836 284
rect 4972 276 4980 284
rect 5084 276 5092 284
rect 5196 276 5204 284
rect 5308 276 5316 284
rect 5452 296 5460 304
rect 5548 296 5556 304
rect 5596 296 5604 304
rect 5644 296 5652 304
rect 5788 296 5796 304
rect 6284 296 6292 304
rect 6460 296 6468 304
rect 6524 294 6532 302
rect 6652 296 6660 304
rect 6716 294 6724 302
rect 6972 296 6980 304
rect 7052 296 7060 304
rect 7068 296 7076 304
rect 7132 296 7140 304
rect 7212 296 7220 304
rect 7260 296 7268 304
rect 7324 294 7332 302
rect 7660 296 7668 304
rect 7740 296 7748 304
rect 7788 296 7796 304
rect 7916 296 7924 304
rect 7980 296 7988 304
rect 8012 296 8020 304
rect 8060 296 8068 304
rect 8092 296 8100 304
rect 5468 276 5476 284
rect 5724 276 5732 284
rect 5788 276 5796 284
rect 5900 276 5908 284
rect 5948 276 5956 284
rect 6108 276 6116 284
rect 6236 276 6244 284
rect 6556 276 6564 284
rect 6812 276 6820 284
rect 6860 276 6868 284
rect 6892 276 6900 284
rect 7036 276 7044 284
rect 7100 276 7108 284
rect 7196 276 7204 284
rect 7228 276 7236 284
rect 7340 276 7348 284
rect 7468 276 7476 284
rect 7708 276 7716 284
rect 7740 276 7748 284
rect 7804 276 7812 284
rect 7820 276 7828 284
rect 7932 276 7940 284
rect 7964 276 7972 284
rect 7996 276 8004 284
rect 8156 276 8164 284
rect 2428 256 2436 264
rect 2620 256 2628 264
rect 2988 256 2996 264
rect 3452 256 3460 264
rect 3740 256 3748 264
rect 3820 256 3828 264
rect 4380 256 4388 264
rect 4572 256 4580 264
rect 4892 256 4900 264
rect 4924 256 4932 264
rect 4956 256 4964 264
rect 5292 256 5300 264
rect 5484 256 5492 264
rect 5548 256 5556 264
rect 5708 256 5716 264
rect 6332 256 6340 264
rect 6796 256 6804 264
rect 6924 256 6932 264
rect 7004 256 7012 264
rect 7260 256 7268 264
rect 7628 256 7636 264
rect 8092 256 8100 264
rect 12 236 20 244
rect 604 236 612 244
rect 844 236 852 244
rect 1308 236 1316 244
rect 1532 236 1540 244
rect 1932 236 1940 244
rect 1948 236 1956 244
rect 2316 236 2324 244
rect 2796 236 2804 244
rect 3388 236 3396 244
rect 4012 236 4020 244
rect 4284 236 4292 244
rect 4796 236 4804 244
rect 5180 236 5188 244
rect 5340 236 5348 244
rect 5852 236 5860 244
rect 6252 236 6260 244
rect 6588 236 6596 244
rect 6780 236 6788 244
rect 6828 236 6836 244
rect 7580 236 7588 244
rect 7692 236 7700 244
rect 7852 236 7860 244
rect 7868 236 7876 244
rect 7948 236 7956 244
rect 8044 236 8052 244
rect 8076 236 8084 244
rect 428 216 436 224
rect 4956 216 4964 224
rect 5548 216 5556 224
rect 3278 206 3286 214
rect 3292 206 3300 214
rect 3306 206 3314 214
rect 6350 206 6358 214
rect 6364 206 6372 214
rect 6378 206 6386 214
rect 5292 196 5300 204
rect 92 176 100 184
rect 204 176 212 184
rect 284 176 292 184
rect 396 176 404 184
rect 556 176 564 184
rect 716 176 724 184
rect 1164 176 1172 184
rect 1196 176 1204 184
rect 1564 176 1572 184
rect 1628 176 1636 184
rect 1692 176 1700 184
rect 1804 176 1812 184
rect 2012 176 2020 184
rect 2172 176 2180 184
rect 2332 176 2340 184
rect 2540 176 2548 184
rect 2748 176 2756 184
rect 2796 176 2804 184
rect 2828 176 2836 184
rect 3036 176 3044 184
rect 3676 176 3684 184
rect 3708 176 3716 184
rect 3820 176 3828 184
rect 3932 176 3940 184
rect 4028 176 4036 184
rect 4300 176 4308 184
rect 4364 176 4372 184
rect 4444 176 4452 184
rect 4492 176 4500 184
rect 4524 176 4532 184
rect 4652 176 4660 184
rect 4940 176 4948 184
rect 5372 176 5380 184
rect 5580 176 5588 184
rect 5772 176 5780 184
rect 7116 176 7124 184
rect 7836 176 7844 184
rect 8092 176 8100 184
rect 76 156 84 164
rect 12 136 20 144
rect 156 136 164 144
rect 460 156 468 164
rect 476 156 484 164
rect 812 156 820 164
rect 1516 156 1524 164
rect 1612 156 1620 164
rect 1644 156 1652 164
rect 1708 156 1716 164
rect 1852 156 1860 164
rect 2188 156 2196 164
rect 2460 156 2468 164
rect 2572 156 2580 164
rect 2764 156 2772 164
rect 2780 156 2788 164
rect 3164 156 3172 164
rect 3228 156 3236 164
rect 3244 156 3252 164
rect 3420 156 3428 164
rect 3532 156 3540 164
rect 3692 156 3700 164
rect 3724 156 3732 164
rect 3772 156 3780 164
rect 3948 156 3956 164
rect 4172 156 4180 164
rect 4316 156 4324 164
rect 4332 156 4340 164
rect 4460 156 4468 164
rect 4540 156 4548 164
rect 4556 156 4564 164
rect 4844 156 4852 164
rect 4924 156 4932 164
rect 5132 156 5140 164
rect 5212 156 5220 164
rect 5228 156 5236 164
rect 5292 156 5300 164
rect 5308 156 5316 164
rect 5564 156 5572 164
rect 5756 156 5764 164
rect 6524 156 6532 164
rect 6668 156 6676 164
rect 6732 156 6740 164
rect 6844 156 6852 164
rect 252 136 260 144
rect 316 136 324 144
rect 412 136 420 144
rect 492 136 500 144
rect 588 136 596 144
rect 668 136 676 144
rect 716 136 724 144
rect 748 136 756 144
rect 828 136 836 144
rect 844 136 852 144
rect 892 136 900 144
rect 940 136 948 144
rect 1148 136 1156 144
rect 1180 136 1188 144
rect 1356 136 1364 144
rect 1388 136 1396 144
rect 1500 136 1508 144
rect 1676 136 1684 144
rect 1724 136 1732 144
rect 1868 136 1876 144
rect 1964 136 1972 144
rect 1996 136 2004 144
rect 2028 136 2036 144
rect 2076 136 2084 144
rect 2108 136 2116 144
rect 2156 136 2164 144
rect 2236 132 2244 140
rect 2252 136 2260 144
rect 2316 136 2324 144
rect 2524 136 2532 144
rect 2604 136 2612 144
rect 2636 136 2644 144
rect 2732 136 2740 144
rect 2844 136 2852 144
rect 2892 136 2900 144
rect 2908 136 2916 144
rect 2988 136 2996 144
rect 3020 136 3028 144
rect 3308 136 3316 144
rect 3404 136 3412 144
rect 3436 136 3444 144
rect 3452 136 3460 144
rect 3740 136 3748 144
rect 3788 136 3796 144
rect 3852 136 3860 144
rect 3884 136 3892 144
rect 7372 156 7380 164
rect 7532 156 7540 164
rect 7852 156 7860 164
rect 4044 136 4052 144
rect 4076 136 4084 144
rect 4108 136 4116 144
rect 4348 136 4356 144
rect 4428 136 4436 144
rect 4508 136 4516 144
rect 4572 136 4580 144
rect 4588 136 4596 144
rect 4700 136 4708 144
rect 4748 136 4756 144
rect 4764 136 4772 144
rect 4860 136 4868 144
rect 5100 136 5108 144
rect 5164 136 5172 144
rect 5260 136 5268 144
rect 5324 136 5332 144
rect 5340 136 5348 144
rect 5532 136 5540 144
rect 5596 136 5604 144
rect 5692 136 5700 144
rect 5724 136 5732 144
rect 5932 136 5940 144
rect 6108 136 6116 144
rect 6236 136 6244 144
rect 6460 136 6468 144
rect 6476 132 6484 140
rect 6588 136 6596 144
rect 6620 136 6628 144
rect 6636 136 6644 144
rect 6716 136 6724 144
rect 6780 136 6788 144
rect 6812 136 6820 144
rect 6844 136 6852 144
rect 6876 136 6884 144
rect 6988 136 6996 144
rect 7276 136 7284 144
rect 7308 136 7316 144
rect 7404 136 7412 144
rect 7580 136 7588 144
rect 7868 136 7876 144
rect 7884 136 7892 144
rect 7932 136 7940 144
rect 7964 136 7972 144
rect 8012 136 8020 144
rect 8044 136 8052 144
rect 28 116 36 124
rect 60 116 68 124
rect 140 116 148 124
rect 236 116 244 124
rect 348 116 356 124
rect 428 116 436 124
rect 444 116 452 124
rect 620 116 628 124
rect 652 116 660 124
rect 668 116 676 124
rect 732 116 740 124
rect 764 116 772 124
rect 1036 116 1044 124
rect 1052 116 1060 124
rect 1260 116 1268 124
rect 1324 118 1332 126
rect 1388 116 1396 124
rect 1420 116 1428 124
rect 1516 116 1524 124
rect 1580 116 1588 124
rect 1820 116 1828 124
rect 1868 116 1876 124
rect 1980 116 1988 124
rect 2044 116 2052 124
rect 2188 116 2196 124
rect 2300 116 2308 124
rect 2460 118 2468 126
rect 2620 116 2628 124
rect 2908 116 2916 124
rect 2924 116 2932 124
rect 188 96 196 104
rect 204 96 212 104
rect 300 96 308 104
rect 348 96 356 104
rect 796 96 804 104
rect 876 96 884 104
rect 940 96 948 104
rect 1148 96 1156 104
rect 1452 96 1460 104
rect 1612 96 1620 104
rect 1756 96 1764 104
rect 1836 96 1844 104
rect 1916 96 1924 104
rect 1932 96 1940 104
rect 2060 96 2068 104
rect 2124 96 2132 104
rect 2252 96 2260 104
rect 2556 96 2564 104
rect 2572 96 2580 104
rect 2668 96 2676 104
rect 2812 96 2820 104
rect 2844 96 2852 104
rect 2956 96 2964 104
rect 3004 116 3012 124
rect 3132 116 3140 124
rect 3340 116 3348 124
rect 3468 116 3476 124
rect 3532 118 3540 126
rect 3836 116 3844 124
rect 3868 116 3876 124
rect 3900 116 3908 124
rect 3916 116 3924 124
rect 3692 96 3700 104
rect 3772 96 3780 104
rect 3820 96 3828 104
rect 3996 96 4004 104
rect 4092 116 4100 124
rect 4172 118 4180 126
rect 4060 96 4068 104
rect 4604 116 4612 124
rect 4396 96 4404 104
rect 4476 96 4484 104
rect 4636 96 4644 104
rect 4684 116 4692 124
rect 4876 116 4884 124
rect 5052 116 5060 124
rect 5180 116 5188 124
rect 5356 116 5364 124
rect 5468 116 5476 124
rect 5708 116 5716 124
rect 5884 116 5892 124
rect 5964 116 5972 124
rect 5980 116 5988 124
rect 6092 116 6100 124
rect 6284 116 6292 124
rect 6524 116 6532 124
rect 6572 116 6580 124
rect 6764 116 6772 124
rect 6796 116 6804 124
rect 6828 116 6836 124
rect 6892 116 6900 124
rect 6940 116 6948 124
rect 6972 116 6980 124
rect 7004 116 7012 124
rect 7052 116 7060 124
rect 7228 116 7236 124
rect 7420 116 7428 124
rect 7596 118 7604 126
rect 7708 118 7716 126
rect 7932 116 7940 124
rect 7948 116 7956 124
rect 7996 116 8004 124
rect 8060 116 8068 124
rect 8092 116 8100 124
rect 4812 96 4820 104
rect 4924 96 4932 104
rect 5148 96 5156 104
rect 5212 96 5220 104
rect 5756 96 5764 104
rect 6012 96 6020 104
rect 6604 96 6612 104
rect 6652 96 6660 104
rect 6668 96 6676 104
rect 6748 96 6756 104
rect 6924 96 6932 104
rect 7020 96 7028 104
rect 7052 96 7060 104
rect 7356 96 7364 104
rect 7388 96 7396 104
rect 7420 96 7428 104
rect 7916 96 7924 104
rect 7980 96 7988 104
rect 8012 96 8020 104
rect 8076 96 8084 104
rect 140 76 148 84
rect 764 76 772 84
rect 956 76 964 84
rect 1532 76 1540 84
rect 1564 76 1572 84
rect 1884 76 1892 84
rect 1964 76 1972 84
rect 3660 76 3668 84
rect 5660 76 5668 84
rect 6204 76 6212 84
rect 6396 76 6404 84
rect 8108 76 8116 84
rect 1742 6 1750 14
rect 1756 6 1764 14
rect 1770 6 1778 14
rect 4814 6 4822 14
rect 4828 6 4836 14
rect 4842 6 4850 14
<< metal2 >>
rect 2365 5764 2371 5776
rect 285 5744 291 5756
rect 125 5704 131 5716
rect 77 5504 83 5576
rect 125 5504 131 5696
rect 205 5664 211 5696
rect 365 5684 371 5736
rect 189 5503 195 5636
rect 301 5524 307 5636
rect 365 5584 371 5656
rect 397 5564 403 5696
rect 429 5684 435 5756
rect 637 5744 643 5756
rect 557 5704 563 5716
rect 637 5684 643 5736
rect 685 5724 691 5756
rect 189 5497 204 5503
rect 125 5344 131 5496
rect 253 5484 259 5516
rect 333 5504 339 5516
rect 189 5444 195 5456
rect 269 5444 275 5496
rect 205 5364 211 5376
rect 125 5104 131 5336
rect 205 5184 211 5356
rect 237 5304 243 5436
rect 285 5383 291 5496
rect 285 5377 300 5383
rect 301 5324 307 5376
rect 317 5364 323 5456
rect 349 5344 355 5476
rect 365 5383 371 5496
rect 397 5464 403 5516
rect 413 5484 419 5636
rect 445 5464 451 5556
rect 477 5484 483 5516
rect 365 5377 387 5383
rect 317 5304 323 5316
rect 349 5304 355 5336
rect 365 5324 371 5356
rect 381 5304 387 5377
rect 413 5344 419 5396
rect 429 5384 435 5456
rect 445 5324 451 5456
rect 461 5364 467 5436
rect 461 5344 467 5356
rect 461 5304 467 5316
rect 429 5284 435 5296
rect 477 5283 483 5336
rect 493 5304 499 5536
rect 541 5524 547 5676
rect 717 5664 723 5696
rect 749 5644 755 5696
rect 909 5684 915 5696
rect 557 5524 563 5556
rect 509 5504 515 5516
rect 541 5404 547 5516
rect 573 5504 579 5536
rect 749 5504 755 5636
rect 909 5604 915 5676
rect 957 5584 963 5596
rect 973 5524 979 5736
rect 989 5724 995 5756
rect 541 5344 547 5396
rect 557 5384 563 5496
rect 573 5384 579 5496
rect 605 5424 611 5456
rect 557 5364 563 5376
rect 621 5364 627 5436
rect 557 5324 563 5356
rect 669 5343 675 5456
rect 653 5337 675 5343
rect 525 5284 531 5296
rect 468 5277 483 5283
rect 237 5084 243 5096
rect 13 4944 19 4956
rect 125 4944 131 5056
rect 77 4904 83 4916
rect 93 4884 99 4936
rect 141 4904 147 4976
rect 189 4924 195 4956
rect 205 4944 211 4996
rect 253 4964 259 5096
rect 269 5043 275 5076
rect 445 5064 451 5256
rect 461 5184 467 5276
rect 541 5144 547 5316
rect 653 5264 659 5337
rect 685 5324 691 5436
rect 701 5344 707 5356
rect 765 5304 771 5476
rect 797 5384 803 5496
rect 989 5484 995 5556
rect 845 5424 851 5476
rect 877 5444 883 5476
rect 893 5464 899 5480
rect 1005 5483 1011 5636
rect 1021 5584 1027 5656
rect 1069 5544 1075 5756
rect 1869 5744 1875 5756
rect 1149 5703 1155 5736
rect 1229 5717 1244 5723
rect 1140 5697 1155 5703
rect 1149 5683 1155 5697
rect 1149 5677 1171 5683
rect 1101 5524 1107 5536
rect 1005 5477 1020 5483
rect 1037 5444 1043 5496
rect 1053 5464 1059 5476
rect 925 5384 931 5436
rect 813 5324 819 5336
rect 829 5324 835 5376
rect 845 5344 851 5376
rect 941 5344 947 5356
rect 973 5344 979 5416
rect 1021 5324 1027 5416
rect 1101 5384 1107 5516
rect 1165 5464 1171 5677
rect 1181 5544 1187 5676
rect 1181 5504 1187 5536
rect 1229 5524 1235 5717
rect 1133 5384 1139 5456
rect 1197 5384 1203 5476
rect 1229 5464 1235 5476
rect 1213 5424 1219 5436
rect 1261 5404 1267 5736
rect 1325 5724 1331 5736
rect 1485 5724 1491 5736
rect 1341 5664 1347 5716
rect 1357 5684 1363 5696
rect 1341 5484 1347 5516
rect 1373 5504 1379 5536
rect 605 5104 611 5216
rect 669 5144 675 5276
rect 269 5037 291 5043
rect 285 5004 291 5037
rect 381 5024 387 5056
rect 285 4944 291 4996
rect 397 4984 403 5036
rect 285 4924 291 4936
rect 173 4904 179 4916
rect 157 4884 163 4896
rect 173 4684 179 4776
rect 189 4744 195 4916
rect 269 4724 275 4916
rect 317 4904 323 4956
rect 365 4924 371 4936
rect 397 4923 403 4976
rect 381 4917 403 4923
rect 381 4904 387 4917
rect 349 4884 355 4896
rect 308 4857 323 4863
rect 285 4724 291 4756
rect 301 4744 307 4836
rect 301 4704 307 4736
rect 173 4544 179 4676
rect 205 4644 211 4656
rect 221 4524 227 4676
rect 253 4664 259 4696
rect 317 4684 323 4857
rect 365 4744 371 4836
rect 381 4784 387 4876
rect 413 4844 419 4916
rect 429 4884 435 4956
rect 445 4824 451 5056
rect 461 5004 467 5036
rect 461 4924 467 4956
rect 461 4904 467 4916
rect 349 4684 355 4716
rect 461 4702 467 4736
rect 477 4724 483 4836
rect 397 4664 403 4696
rect 253 4584 259 4636
rect 13 4404 19 4436
rect 68 4297 83 4303
rect 13 3984 19 4136
rect 29 4124 35 4236
rect 77 4184 83 4297
rect 93 4284 99 4516
rect 109 4324 115 4396
rect 109 4243 115 4316
rect 141 4304 147 4356
rect 173 4304 179 4316
rect 109 4237 131 4243
rect 109 4144 115 4216
rect 125 4124 131 4237
rect 173 4144 179 4156
rect 189 4144 195 4236
rect 205 4204 211 4516
rect 237 4344 243 4516
rect 301 4504 307 4516
rect 317 4504 323 4576
rect 349 4564 355 4576
rect 388 4517 403 4523
rect 381 4504 387 4516
rect 285 4497 300 4503
rect 237 4284 243 4336
rect 253 4264 259 4436
rect 285 4324 291 4497
rect 301 4364 307 4476
rect 397 4384 403 4517
rect 429 4483 435 4536
rect 477 4504 483 4536
rect 413 4477 435 4483
rect 301 4324 307 4356
rect 285 4304 291 4316
rect 349 4304 355 4356
rect 349 4284 355 4296
rect 381 4284 387 4316
rect 413 4284 419 4477
rect 477 4284 483 4296
rect 205 4164 211 4176
rect 237 4140 243 4256
rect 333 4224 339 4276
rect 413 4264 419 4276
rect 493 4264 499 5096
rect 813 5084 819 5296
rect 909 5184 915 5316
rect 1133 5304 1139 5376
rect 1149 5344 1155 5376
rect 1213 5350 1219 5396
rect 1277 5384 1283 5480
rect 1293 5464 1299 5476
rect 1293 5344 1299 5456
rect 1309 5404 1315 5476
rect 1309 5364 1315 5376
rect 1245 5324 1251 5336
rect 1293 5324 1299 5336
rect 1117 5104 1123 5136
rect 1181 5124 1187 5196
rect 1309 5164 1315 5356
rect 1357 5304 1363 5316
rect 1389 5304 1395 5476
rect 1405 5444 1411 5516
rect 1421 5484 1427 5696
rect 1581 5684 1587 5696
rect 1469 5544 1475 5676
rect 1405 5384 1411 5436
rect 1485 5424 1491 5456
rect 1517 5344 1523 5676
rect 1565 5544 1571 5636
rect 1597 5584 1603 5716
rect 1645 5704 1651 5716
rect 1613 5664 1619 5696
rect 1629 5564 1635 5696
rect 1613 5502 1619 5536
rect 1661 5504 1667 5736
rect 1677 5704 1683 5716
rect 1597 5364 1603 5396
rect 1645 5384 1651 5456
rect 1645 5364 1651 5376
rect 1277 5124 1283 5136
rect 1357 5124 1363 5196
rect 525 5044 531 5056
rect 509 4924 515 5036
rect 509 4884 515 4916
rect 525 4884 531 5036
rect 557 4944 563 4956
rect 557 4904 563 4916
rect 557 4864 563 4876
rect 525 4704 531 4776
rect 509 4524 515 4536
rect 525 4524 531 4556
rect 557 4503 563 4516
rect 548 4497 563 4503
rect 573 4304 579 5076
rect 637 4984 643 5076
rect 685 4944 691 5076
rect 589 4884 595 4896
rect 653 4884 659 4936
rect 589 4704 595 4736
rect 605 4644 611 4716
rect 621 4644 627 4816
rect 685 4784 691 4936
rect 717 4904 723 4918
rect 701 4704 707 4836
rect 637 4684 643 4696
rect 717 4684 723 4776
rect 749 4704 755 4856
rect 621 4564 627 4636
rect 589 4324 595 4436
rect 253 4144 259 4216
rect 365 4204 371 4236
rect 29 3904 35 4036
rect 77 4024 83 4096
rect 237 3904 243 4132
rect 29 3844 35 3856
rect 125 3744 131 3876
rect 205 3764 211 3896
rect 253 3883 259 4136
rect 269 4104 275 4196
rect 429 4124 435 4176
rect 317 4024 323 4036
rect 445 4024 451 4256
rect 525 4243 531 4276
rect 509 4237 531 4243
rect 493 4184 499 4236
rect 509 4224 515 4237
rect 509 4184 515 4216
rect 541 4124 547 4236
rect 557 4164 563 4196
rect 621 4164 627 4556
rect 717 4544 723 4676
rect 733 4664 739 4696
rect 781 4584 787 4976
rect 813 4944 819 5076
rect 829 4964 835 5036
rect 813 4704 819 4736
rect 829 4724 835 4956
rect 877 4924 883 5096
rect 973 4984 979 5056
rect 1069 4984 1075 5076
rect 1117 4984 1123 5056
rect 1005 4944 1011 4956
rect 1149 4924 1155 4996
rect 1181 4964 1187 5036
rect 1213 4984 1219 5096
rect 1229 5044 1235 5076
rect 1245 5064 1251 5076
rect 1261 4984 1267 5036
rect 893 4784 899 4876
rect 973 4724 979 4836
rect 829 4683 835 4696
rect 820 4677 835 4683
rect 877 4684 883 4716
rect 861 4624 867 4680
rect 909 4624 915 4656
rect 973 4604 979 4694
rect 1133 4664 1139 4716
rect 1181 4684 1187 4956
rect 1197 4944 1203 4956
rect 1229 4904 1235 4936
rect 1277 4923 1283 5116
rect 1309 5084 1315 5096
rect 1309 4944 1315 5056
rect 1309 4924 1315 4936
rect 1325 4924 1331 5096
rect 1341 5064 1347 5116
rect 1389 5083 1395 5136
rect 1517 5104 1523 5336
rect 1613 5204 1619 5236
rect 1661 5102 1667 5396
rect 1677 5384 1683 5696
rect 1693 5684 1699 5736
rect 1789 5664 1795 5696
rect 1837 5644 1843 5736
rect 1736 5606 1742 5614
rect 1750 5606 1756 5614
rect 1764 5606 1770 5614
rect 1778 5606 1784 5614
rect 1821 5463 1827 5636
rect 1885 5584 1891 5636
rect 1853 5504 1859 5536
rect 1812 5457 1827 5463
rect 1757 5444 1763 5456
rect 1677 5344 1683 5376
rect 1709 5224 1715 5316
rect 1757 5284 1763 5436
rect 1736 5206 1742 5214
rect 1750 5206 1756 5214
rect 1764 5206 1770 5214
rect 1778 5206 1784 5214
rect 1805 5184 1811 5416
rect 1821 5404 1827 5436
rect 1837 5384 1843 5476
rect 1901 5444 1907 5676
rect 1981 5664 1987 5736
rect 2173 5544 2179 5636
rect 2253 5584 2259 5716
rect 1949 5517 1964 5523
rect 1949 5484 1955 5517
rect 1901 5344 1907 5436
rect 1949 5384 1955 5476
rect 1965 5364 1971 5436
rect 1981 5384 1987 5496
rect 2029 5464 2035 5516
rect 2093 5504 2099 5536
rect 2157 5504 2163 5536
rect 2173 5503 2179 5536
rect 2221 5524 2227 5536
rect 2173 5497 2195 5503
rect 1981 5324 1987 5376
rect 1997 5364 2003 5456
rect 2029 5424 2035 5456
rect 2045 5384 2051 5396
rect 1997 5284 2003 5356
rect 1917 5104 1923 5116
rect 2029 5104 2035 5136
rect 1469 5084 1475 5094
rect 1517 5084 1523 5096
rect 1373 5077 1395 5083
rect 1268 4917 1283 4923
rect 1325 4884 1331 4916
rect 1357 4904 1363 5036
rect 1373 4984 1379 5077
rect 1421 4944 1427 4956
rect 1261 4724 1267 4836
rect 1293 4784 1299 4876
rect 1357 4864 1363 4896
rect 1261 4664 1267 4696
rect 1309 4684 1315 4756
rect 1117 4644 1123 4656
rect 861 4584 867 4596
rect 1101 4584 1107 4636
rect 685 4324 691 4496
rect 701 4324 707 4336
rect 637 4284 643 4296
rect 685 4284 691 4316
rect 717 4144 723 4536
rect 781 4364 787 4576
rect 1005 4564 1011 4576
rect 1133 4564 1139 4656
rect 852 4537 867 4543
rect 861 4384 867 4537
rect 781 4303 787 4356
rect 765 4297 787 4303
rect 765 4264 771 4297
rect 813 4264 819 4296
rect 893 4144 899 4156
rect 925 4144 931 4396
rect 941 4344 947 4516
rect 957 4404 963 4556
rect 973 4343 979 4436
rect 989 4364 995 4516
rect 973 4337 995 4343
rect 989 4324 995 4337
rect 973 4304 979 4316
rect 941 4144 947 4276
rect 1005 4184 1011 4556
rect 1037 4464 1043 4516
rect 1165 4504 1171 4636
rect 1181 4624 1187 4656
rect 1293 4540 1299 4676
rect 1085 4384 1091 4476
rect 1133 4384 1139 4456
rect 1245 4437 1260 4443
rect 1149 4344 1155 4356
rect 1053 4284 1059 4296
rect 1037 4264 1043 4276
rect 1005 4144 1011 4176
rect 1053 4164 1059 4276
rect 541 4064 547 4116
rect 589 4044 595 4096
rect 653 4063 659 4116
rect 676 4077 691 4083
rect 653 4057 675 4063
rect 477 3944 483 4016
rect 244 3877 259 3883
rect 125 3724 131 3736
rect 93 3584 99 3716
rect 45 3464 51 3496
rect 13 3364 19 3436
rect 93 3384 99 3496
rect 109 3444 115 3536
rect 157 3464 163 3696
rect 221 3504 227 3836
rect 253 3724 259 3836
rect 413 3724 419 3856
rect 493 3724 499 3736
rect 269 3704 275 3716
rect 285 3704 291 3716
rect 349 3704 355 3718
rect 413 3604 419 3716
rect 461 3504 467 3696
rect 477 3484 483 3636
rect 141 3384 147 3456
rect 45 3284 51 3336
rect 61 3283 67 3316
rect 77 3304 83 3336
rect 61 3277 76 3283
rect 13 3103 19 3236
rect 61 3144 67 3277
rect 93 3124 99 3316
rect 13 3097 35 3103
rect 13 3064 19 3076
rect 13 2944 19 3056
rect 29 2944 35 3097
rect 45 2944 51 3116
rect 93 3104 99 3116
rect 141 3104 147 3296
rect 157 3104 163 3456
rect 173 3424 179 3456
rect 237 3384 243 3436
rect 253 3424 259 3456
rect 141 3084 147 3096
rect 157 3084 163 3096
rect 173 3084 179 3336
rect 189 3324 195 3336
rect 205 3304 211 3316
rect 237 3304 243 3356
rect 349 3324 355 3336
rect 349 3283 355 3316
rect 381 3303 387 3476
rect 477 3464 483 3476
rect 509 3444 515 3876
rect 525 3864 531 3896
rect 541 3884 547 3956
rect 525 3724 531 3856
rect 573 3764 579 3936
rect 589 3924 595 4036
rect 669 3984 675 4057
rect 685 4044 691 4077
rect 733 3984 739 4036
rect 589 3764 595 3816
rect 621 3784 627 3896
rect 637 3884 643 3916
rect 653 3823 659 3916
rect 685 3864 691 3936
rect 653 3817 668 3823
rect 669 3744 675 3816
rect 685 3703 691 3856
rect 717 3744 723 3876
rect 733 3744 739 3896
rect 765 3744 771 3776
rect 701 3724 707 3736
rect 781 3724 787 3896
rect 829 3824 835 3876
rect 685 3697 700 3703
rect 797 3624 803 3736
rect 845 3724 851 3896
rect 861 3864 867 4136
rect 925 4044 931 4136
rect 957 4104 963 4136
rect 1021 4044 1027 4156
rect 1053 4124 1059 4156
rect 1101 4144 1107 4276
rect 1117 4264 1123 4316
rect 1245 4304 1251 4437
rect 1261 4324 1267 4356
rect 1252 4297 1267 4303
rect 1133 4284 1139 4296
rect 1181 4284 1187 4296
rect 1229 4284 1235 4296
rect 1069 4104 1075 4116
rect 1085 4084 1091 4136
rect 1117 4124 1123 4136
rect 1133 4124 1139 4196
rect 1197 4124 1203 4236
rect 1245 4164 1251 4176
rect 1053 3884 1059 3916
rect 893 3864 899 3876
rect 861 3804 867 3856
rect 909 3824 915 3876
rect 1021 3864 1027 3876
rect 893 3764 899 3796
rect 813 3664 819 3716
rect 861 3703 867 3736
rect 893 3724 899 3756
rect 925 3744 931 3756
rect 973 3724 979 3776
rect 1021 3740 1027 3756
rect 1037 3744 1043 3816
rect 989 3724 995 3736
rect 1053 3724 1059 3876
rect 1069 3784 1075 3836
rect 1085 3744 1091 4036
rect 1101 3884 1107 3936
rect 1149 3904 1155 4056
rect 1165 3984 1171 4076
rect 1261 4044 1267 4297
rect 1277 3923 1283 4516
rect 1293 4264 1299 4276
rect 1277 3917 1299 3923
rect 1213 3884 1219 3916
rect 1117 3744 1123 3836
rect 852 3697 867 3703
rect 909 3684 915 3716
rect 1101 3684 1107 3736
rect 1117 3704 1123 3716
rect 477 3437 492 3443
rect 397 3384 403 3436
rect 461 3304 467 3336
rect 381 3297 396 3303
rect 333 3277 355 3283
rect 333 3144 339 3277
rect 333 3123 339 3136
rect 381 3124 387 3236
rect 324 3117 339 3123
rect 237 3104 243 3116
rect 93 2964 99 3036
rect 45 2924 51 2936
rect 45 2864 51 2896
rect 61 2702 67 2936
rect 77 2864 83 2956
rect 109 2684 115 3036
rect 141 2944 147 3076
rect 173 3064 179 3076
rect 189 3044 195 3080
rect 221 2944 227 3036
rect 253 2944 259 3036
rect 141 2904 147 2916
rect 157 2724 163 2916
rect 317 2903 323 3036
rect 365 2964 371 3096
rect 429 3084 435 3296
rect 477 3144 483 3437
rect 525 3424 531 3496
rect 573 3484 579 3596
rect 813 3504 819 3636
rect 941 3584 947 3616
rect 493 3384 499 3416
rect 509 3304 515 3396
rect 525 3284 531 3316
rect 541 3284 547 3316
rect 589 3304 595 3316
rect 525 3084 531 3156
rect 429 3044 435 3076
rect 541 3064 547 3136
rect 557 3064 563 3236
rect 605 3184 611 3216
rect 621 3204 627 3496
rect 637 3344 643 3476
rect 973 3464 979 3676
rect 1005 3504 1011 3536
rect 957 3444 963 3456
rect 733 3404 739 3436
rect 637 3304 643 3336
rect 685 3324 691 3336
rect 669 3264 675 3316
rect 637 3124 643 3176
rect 685 3163 691 3316
rect 676 3157 691 3163
rect 621 3117 636 3123
rect 573 3084 579 3116
rect 621 3064 627 3117
rect 669 3084 675 3156
rect 701 3144 707 3256
rect 717 3244 723 3356
rect 733 3304 739 3316
rect 749 3264 755 3316
rect 765 3284 771 3316
rect 797 3284 803 3396
rect 989 3363 995 3436
rect 989 3357 1011 3363
rect 1005 3344 1011 3357
rect 989 3324 995 3336
rect 733 3184 739 3196
rect 733 3084 739 3096
rect 717 3064 723 3076
rect 317 2897 332 2903
rect 189 2784 195 2856
rect 237 2784 243 2876
rect 365 2864 371 2936
rect 461 2924 467 2996
rect 269 2744 275 2836
rect 397 2724 403 2736
rect 317 2704 323 2716
rect 29 2584 35 2676
rect 269 2544 275 2696
rect 429 2684 435 2696
rect 477 2684 483 3064
rect 557 3004 563 3036
rect 621 2984 627 3056
rect 493 2924 499 2936
rect 637 2924 643 3056
rect 685 3044 691 3056
rect 493 2704 499 2916
rect 749 2884 755 3236
rect 765 3224 771 3276
rect 781 3104 787 3136
rect 797 3103 803 3276
rect 829 3124 835 3236
rect 925 3224 931 3296
rect 941 3264 947 3316
rect 1005 3244 1011 3316
rect 1021 3304 1027 3496
rect 1037 3364 1043 3676
rect 1133 3524 1139 3576
rect 1053 3504 1059 3516
rect 1117 3464 1123 3476
rect 1149 3384 1155 3876
rect 1197 3864 1203 3880
rect 1197 3744 1203 3856
rect 1245 3844 1251 3856
rect 1261 3844 1267 3876
rect 1277 3764 1283 3896
rect 1293 3804 1299 3917
rect 1309 3884 1315 4676
rect 1325 4664 1331 4694
rect 1421 4604 1427 4936
rect 1453 4924 1459 4956
rect 1485 4923 1491 4956
rect 1549 4944 1555 4976
rect 1485 4917 1500 4923
rect 1453 4804 1459 4916
rect 1517 4904 1523 4936
rect 1597 4923 1603 5036
rect 1588 4917 1603 4923
rect 1437 4684 1443 4736
rect 1485 4724 1491 4796
rect 1549 4743 1555 4836
rect 1549 4737 1571 4743
rect 1453 4684 1459 4716
rect 1485 4684 1491 4716
rect 1549 4604 1555 4716
rect 1325 4584 1331 4596
rect 1533 4544 1539 4556
rect 1357 4304 1363 4356
rect 1373 4164 1379 4476
rect 1389 4344 1395 4436
rect 1469 4384 1475 4518
rect 1501 4504 1507 4536
rect 1565 4523 1571 4737
rect 1581 4684 1587 4916
rect 1597 4844 1603 4876
rect 1597 4704 1603 4836
rect 1629 4764 1635 5076
rect 2045 5064 2051 5376
rect 2061 5344 2067 5436
rect 2109 5343 2115 5476
rect 2125 5344 2131 5476
rect 2100 5337 2115 5343
rect 2141 5324 2147 5456
rect 2173 5344 2179 5376
rect 2189 5324 2195 5497
rect 2205 5344 2211 5356
rect 2285 5344 2291 5716
rect 2333 5584 2339 5696
rect 2413 5684 2419 5716
rect 2077 5304 2083 5316
rect 2109 5284 2115 5316
rect 2141 5184 2147 5316
rect 2221 5264 2227 5316
rect 2269 5284 2275 5336
rect 2301 5304 2307 5436
rect 2317 5424 2323 5456
rect 2349 5344 2355 5516
rect 2429 5504 2435 5843
rect 2509 5744 2515 5843
rect 2605 5837 2627 5843
rect 2477 5684 2483 5696
rect 2541 5664 2547 5736
rect 2573 5724 2579 5736
rect 2589 5724 2595 5756
rect 2605 5744 2611 5837
rect 2813 5804 2819 5843
rect 3069 5804 3075 5843
rect 3272 5806 3278 5814
rect 3286 5806 3292 5814
rect 3300 5806 3306 5814
rect 3314 5806 3320 5814
rect 3613 5804 3619 5843
rect 2733 5764 2739 5776
rect 2653 5724 2659 5736
rect 2637 5684 2643 5696
rect 2445 5584 2451 5656
rect 2541 5524 2547 5636
rect 2637 5524 2643 5676
rect 2669 5664 2675 5736
rect 2701 5724 2707 5736
rect 2733 5724 2739 5756
rect 2669 5544 2675 5636
rect 2701 5584 2707 5716
rect 2781 5684 2787 5716
rect 2717 5504 2723 5676
rect 2669 5484 2675 5496
rect 2381 5404 2387 5456
rect 2413 5344 2419 5356
rect 2605 5344 2611 5436
rect 2349 5184 2355 5336
rect 2397 5304 2403 5316
rect 2365 5264 2371 5296
rect 2637 5284 2643 5356
rect 2701 5326 2707 5476
rect 2765 5464 2771 5496
rect 2797 5484 2803 5576
rect 2829 5484 2835 5656
rect 2845 5504 2851 5796
rect 3021 5744 3027 5796
rect 3069 5724 3075 5796
rect 3149 5764 3155 5776
rect 3053 5684 3059 5696
rect 3085 5664 3091 5736
rect 3085 5604 3091 5636
rect 3117 5584 3123 5736
rect 3149 5724 3155 5756
rect 3357 5724 3363 5736
rect 3453 5724 3459 5736
rect 3549 5724 3555 5736
rect 3197 5684 3203 5716
rect 2909 5524 2915 5536
rect 3149 5524 3155 5596
rect 3357 5504 3363 5716
rect 3533 5684 3539 5696
rect 3533 5524 3539 5676
rect 3629 5664 3635 5676
rect 3533 5504 3539 5516
rect 3565 5484 3571 5496
rect 3581 5484 3587 5496
rect 3597 5484 3603 5576
rect 3629 5484 3635 5656
rect 3645 5504 3651 5796
rect 3668 5777 3683 5783
rect 3677 5764 3683 5777
rect 3805 5744 3811 5843
rect 3917 5837 3939 5843
rect 3933 5784 3939 5837
rect 3677 5484 3683 5716
rect 3725 5704 3731 5716
rect 3837 5684 3843 5736
rect 3885 5724 3891 5756
rect 3949 5724 3955 5756
rect 4029 5744 4035 5843
rect 4157 5777 4172 5783
rect 4157 5764 4163 5777
rect 4381 5764 4387 5843
rect 6205 5804 6211 5843
rect 6344 5806 6350 5814
rect 6358 5806 6364 5814
rect 6372 5806 6378 5814
rect 6386 5806 6392 5814
rect 2941 5464 2947 5476
rect 2765 5404 2771 5456
rect 2829 5423 2835 5436
rect 2829 5417 2851 5423
rect 2829 5384 2835 5396
rect 2845 5384 2851 5417
rect 2861 5324 2867 5436
rect 3005 5344 3011 5456
rect 3037 5384 3043 5476
rect 3101 5384 3107 5456
rect 3133 5424 3139 5436
rect 3133 5364 3139 5416
rect 3165 5364 3171 5436
rect 3213 5384 3219 5476
rect 3421 5444 3427 5476
rect 3517 5464 3523 5476
rect 3709 5464 3715 5494
rect 3837 5464 3843 5636
rect 3901 5604 3907 5716
rect 3965 5584 3971 5736
rect 3997 5684 4003 5736
rect 4109 5704 4115 5716
rect 4013 5484 4019 5616
rect 4045 5524 4051 5636
rect 4109 5604 4115 5696
rect 4205 5624 4211 5676
rect 4333 5644 4339 5736
rect 4093 5484 4099 5596
rect 4173 5584 4179 5596
rect 4125 5504 4131 5516
rect 4221 5504 4227 5516
rect 4205 5497 4220 5503
rect 3229 5364 3235 5416
rect 3272 5406 3278 5414
rect 3286 5406 3292 5414
rect 3300 5406 3306 5414
rect 3314 5406 3320 5414
rect 3053 5304 3059 5336
rect 3101 5304 3107 5356
rect 2157 5084 2163 5096
rect 2221 5084 2227 5136
rect 2237 5104 2243 5116
rect 2253 5084 2259 5116
rect 2141 5064 2147 5076
rect 2013 4884 2019 4916
rect 1736 4806 1742 4814
rect 1750 4806 1756 4814
rect 1764 4806 1770 4814
rect 1778 4806 1784 4814
rect 1645 4704 1651 4776
rect 1629 4664 1635 4676
rect 1709 4664 1715 4696
rect 1821 4684 1827 4716
rect 1853 4684 1859 4696
rect 1901 4684 1907 4716
rect 1981 4704 1987 4836
rect 2045 4764 2051 5056
rect 2093 4904 2099 5036
rect 2109 5024 2115 5056
rect 2125 4964 2131 4976
rect 2093 4804 2099 4876
rect 2157 4864 2163 4916
rect 2173 4904 2179 5076
rect 2269 4924 2275 5076
rect 2301 5004 2307 5076
rect 2285 4997 2300 5003
rect 2285 4944 2291 4997
rect 2397 4944 2403 5076
rect 2429 5064 2435 5096
rect 2445 4944 2451 5056
rect 2301 4924 2307 4936
rect 2237 4904 2243 4916
rect 2253 4884 2259 4916
rect 2333 4904 2339 4916
rect 2365 4904 2371 4936
rect 2381 4904 2387 4916
rect 2461 4904 2467 5116
rect 2493 5104 2499 5116
rect 2573 5104 2579 5116
rect 2589 5084 2595 5116
rect 2621 5104 2627 5116
rect 2669 5084 2675 5116
rect 2733 5102 2739 5116
rect 2477 4944 2483 5076
rect 2493 4923 2499 4956
rect 2541 4944 2547 5076
rect 2573 4964 2579 4996
rect 2525 4924 2531 4936
rect 2589 4924 2595 4976
rect 2701 4924 2707 5056
rect 2733 4944 2739 4976
rect 2749 4924 2755 5136
rect 2797 5104 2803 5276
rect 3021 5224 3027 5236
rect 2893 4944 2899 5036
rect 2925 5004 2931 5116
rect 3005 5084 3011 5096
rect 3053 5084 3059 5296
rect 3165 5224 3171 5336
rect 3325 5304 3331 5336
rect 3357 5326 3363 5356
rect 3501 5304 3507 5376
rect 3213 5264 3219 5296
rect 3549 5264 3555 5336
rect 3613 5304 3619 5436
rect 3629 5384 3635 5456
rect 3837 5424 3843 5436
rect 3853 5423 3859 5436
rect 3853 5417 3875 5423
rect 3485 5244 3491 5256
rect 2957 5064 2963 5076
rect 2909 4964 2915 4976
rect 3005 4944 3011 5016
rect 3021 4944 3027 5076
rect 3053 5024 3059 5076
rect 3117 4964 3123 5216
rect 3245 5124 3251 5236
rect 3245 5097 3260 5103
rect 3213 5004 3219 5076
rect 3213 4943 3219 4996
rect 3229 4984 3235 5056
rect 3245 4983 3251 5097
rect 3421 5084 3427 5096
rect 3272 5006 3278 5014
rect 3286 5006 3292 5014
rect 3300 5006 3306 5014
rect 3314 5006 3320 5014
rect 3245 4977 3260 4983
rect 3341 4983 3347 5056
rect 3325 4977 3347 4983
rect 3325 4964 3331 4977
rect 3213 4937 3228 4943
rect 2484 4917 2499 4923
rect 2765 4904 2771 4936
rect 2813 4924 2819 4936
rect 2781 4904 2787 4916
rect 2461 4884 2467 4896
rect 2877 4884 2883 4916
rect 2973 4904 2979 4918
rect 3181 4904 3187 4916
rect 3149 4864 3155 4896
rect 3133 4803 3139 4836
rect 3133 4797 3155 4803
rect 2045 4702 2051 4736
rect 2109 4704 2115 4716
rect 1556 4517 1571 4523
rect 1581 4504 1587 4516
rect 1613 4504 1619 4536
rect 1677 4524 1683 4636
rect 1805 4584 1811 4680
rect 1853 4584 1859 4656
rect 1693 4524 1699 4536
rect 1736 4406 1742 4414
rect 1750 4406 1756 4414
rect 1764 4406 1770 4414
rect 1778 4406 1784 4414
rect 1389 4204 1395 4336
rect 1405 4304 1411 4316
rect 1437 4304 1443 4316
rect 1405 4264 1411 4276
rect 1373 3984 1379 4116
rect 1389 3924 1395 3936
rect 1405 3923 1411 4256
rect 1437 4184 1443 4296
rect 1517 4164 1523 4256
rect 1533 4184 1539 4256
rect 1453 4140 1459 4156
rect 1565 4143 1571 4280
rect 1629 4264 1635 4296
rect 1581 4144 1587 4156
rect 1597 4144 1603 4236
rect 1565 4137 1580 4143
rect 1613 4137 1628 4143
rect 1533 4104 1539 4136
rect 1613 4124 1619 4137
rect 1709 4124 1715 4256
rect 1757 4124 1763 4156
rect 1629 4104 1635 4116
rect 1645 4104 1651 4116
rect 1421 3984 1427 4076
rect 1533 4064 1539 4096
rect 1396 3917 1411 3923
rect 1421 3904 1427 3976
rect 1693 3944 1699 4036
rect 1736 4006 1742 4014
rect 1750 4006 1756 4014
rect 1764 4006 1770 4014
rect 1778 4006 1784 4014
rect 1309 3764 1315 3876
rect 1213 3704 1219 3716
rect 1245 3684 1251 3756
rect 1181 3484 1187 3496
rect 1165 3464 1171 3476
rect 1229 3404 1235 3436
rect 1245 3383 1251 3676
rect 1309 3584 1315 3718
rect 1293 3544 1299 3556
rect 1341 3524 1347 3816
rect 1437 3784 1443 3796
rect 1469 3764 1475 3816
rect 1517 3764 1523 3796
rect 1581 3784 1587 3916
rect 1805 3904 1811 4436
rect 1821 4304 1827 4516
rect 1837 4304 1843 4436
rect 1837 4184 1843 4296
rect 1821 4144 1827 4156
rect 1853 4124 1859 4176
rect 1869 4144 1875 4236
rect 1901 4184 1907 4636
rect 1917 4604 1923 4636
rect 1981 4544 1987 4696
rect 2061 4564 2067 4596
rect 2077 4584 2083 4676
rect 2093 4544 2099 4636
rect 2125 4584 2131 4696
rect 2157 4664 2163 4716
rect 2173 4704 2179 4716
rect 2237 4684 2243 4776
rect 2285 4704 2291 4736
rect 2413 4704 2419 4716
rect 2141 4584 2147 4636
rect 1981 4524 1987 4536
rect 1997 4464 2003 4518
rect 2221 4484 2227 4676
rect 2301 4644 2307 4656
rect 2365 4544 2371 4656
rect 2381 4644 2387 4696
rect 2397 4563 2403 4676
rect 2429 4664 2435 4676
rect 2397 4557 2412 4563
rect 2045 4384 2051 4456
rect 1981 4337 1996 4343
rect 1917 4304 1923 4316
rect 1981 4303 1987 4337
rect 1972 4297 1987 4303
rect 1965 4244 1971 4276
rect 1981 4224 1987 4297
rect 1981 4184 1987 4216
rect 2013 4184 2019 4296
rect 2013 4164 2019 4176
rect 1901 4104 1907 4136
rect 1917 4124 1923 4156
rect 1997 4064 2003 4156
rect 2029 4144 2035 4316
rect 2077 4284 2083 4296
rect 2109 4264 2115 4436
rect 2237 4324 2243 4336
rect 2109 4184 2115 4196
rect 2141 4144 2147 4256
rect 2045 4124 2051 4136
rect 2157 4104 2163 4236
rect 2173 4224 2179 4256
rect 2189 4144 2195 4276
rect 2205 4244 2211 4296
rect 2253 4264 2259 4276
rect 2269 4164 2275 4296
rect 2301 4164 2307 4536
rect 2413 4524 2419 4556
rect 2445 4524 2451 4696
rect 2461 4684 2467 4756
rect 2461 4664 2467 4676
rect 2477 4644 2483 4696
rect 2477 4604 2483 4636
rect 2365 4504 2371 4516
rect 2381 4464 2387 4496
rect 2445 4484 2451 4496
rect 2477 4484 2483 4596
rect 2525 4544 2531 4676
rect 2541 4564 2547 4676
rect 2525 4524 2531 4536
rect 2509 4517 2524 4523
rect 2509 4504 2515 4517
rect 2541 4504 2547 4516
rect 2317 4264 2323 4296
rect 2189 4124 2195 4136
rect 1885 3984 1891 4036
rect 1901 3904 1907 4036
rect 1933 3924 1939 3936
rect 1661 3864 1667 3896
rect 1757 3864 1763 3896
rect 1613 3823 1619 3836
rect 1597 3817 1619 3823
rect 1597 3724 1603 3817
rect 1709 3744 1715 3756
rect 1725 3744 1731 3836
rect 1821 3824 1827 3876
rect 1869 3843 1875 3896
rect 1853 3837 1875 3843
rect 1613 3724 1619 3736
rect 1373 3544 1379 3556
rect 1261 3464 1267 3516
rect 1325 3424 1331 3516
rect 1341 3484 1347 3516
rect 1357 3504 1363 3536
rect 1437 3524 1443 3636
rect 1453 3584 1459 3636
rect 1437 3504 1443 3516
rect 1373 3484 1379 3496
rect 1453 3484 1459 3576
rect 1485 3544 1491 3716
rect 1549 3664 1555 3716
rect 1517 3564 1523 3656
rect 1581 3584 1587 3696
rect 1501 3504 1507 3536
rect 1517 3524 1523 3556
rect 1613 3544 1619 3636
rect 1565 3484 1571 3496
rect 1597 3464 1603 3516
rect 1629 3504 1635 3516
rect 1661 3504 1667 3656
rect 1805 3644 1811 3736
rect 1821 3684 1827 3716
rect 1736 3606 1742 3614
rect 1750 3606 1756 3614
rect 1764 3606 1770 3614
rect 1778 3606 1784 3614
rect 1645 3484 1651 3496
rect 1708 3464 1716 3470
rect 1245 3377 1260 3383
rect 845 3184 851 3196
rect 1021 3184 1027 3296
rect 1037 3284 1043 3316
rect 1101 3304 1107 3336
rect 1069 3204 1075 3296
rect 797 3097 812 3103
rect 893 3084 899 3096
rect 765 2984 771 3056
rect 781 2944 787 2956
rect 797 2944 803 2976
rect 733 2784 739 2836
rect 509 2704 515 2756
rect 749 2744 755 2856
rect 781 2844 787 2936
rect 813 2884 819 3056
rect 829 2984 835 3076
rect 877 3063 883 3076
rect 877 3057 899 3063
rect 829 2784 835 2956
rect 845 2904 851 3036
rect 893 2984 899 3057
rect 957 2944 963 3076
rect 1005 3004 1011 3096
rect 1053 3084 1059 3156
rect 1229 3144 1235 3376
rect 1325 3364 1331 3376
rect 1389 3364 1395 3396
rect 1485 3364 1491 3436
rect 1613 3404 1619 3456
rect 1741 3384 1747 3416
rect 1789 3404 1795 3476
rect 1757 3364 1763 3396
rect 1277 3164 1283 3236
rect 1277 3124 1283 3136
rect 1165 3044 1171 3096
rect 1181 3084 1187 3096
rect 1213 3064 1219 3076
rect 877 2903 883 2936
rect 877 2897 899 2903
rect 845 2784 851 2896
rect 877 2884 883 2897
rect 893 2744 899 2897
rect 605 2702 611 2716
rect 477 2644 483 2656
rect 477 2526 483 2596
rect 509 2564 515 2696
rect 573 2684 579 2696
rect 541 2584 547 2636
rect 285 2443 291 2518
rect 509 2504 515 2536
rect 285 2437 307 2443
rect 29 2284 35 2436
rect 77 2204 83 2296
rect 109 2144 115 2276
rect 157 2224 163 2436
rect 301 2384 307 2437
rect 205 2244 211 2316
rect 221 2244 227 2256
rect 157 2184 163 2196
rect 189 2164 195 2216
rect 13 2084 19 2136
rect 125 2124 131 2136
rect 141 2124 147 2136
rect 173 2124 179 2156
rect 205 2144 211 2236
rect 221 2144 227 2236
rect 237 2204 243 2276
rect 269 2244 275 2316
rect 253 2143 259 2236
rect 285 2223 291 2316
rect 301 2304 307 2356
rect 349 2344 355 2436
rect 324 2337 339 2343
rect 237 2137 259 2143
rect 269 2217 291 2223
rect 29 1784 35 1896
rect 77 1744 83 2076
rect 221 1964 227 2136
rect 237 2124 243 2137
rect 269 2104 275 2217
rect 285 2144 291 2196
rect 253 1984 259 2076
rect 212 1937 227 1943
rect 205 1904 211 1916
rect 221 1904 227 1937
rect 269 1904 275 2096
rect 285 2084 291 2136
rect 301 2124 307 2236
rect 333 2184 339 2337
rect 381 2324 387 2336
rect 349 2284 355 2316
rect 365 2204 371 2296
rect 477 2284 483 2396
rect 509 2304 515 2316
rect 525 2297 540 2303
rect 397 2124 403 2196
rect 413 2144 419 2276
rect 477 2264 483 2276
rect 429 2144 435 2236
rect 461 2144 467 2236
rect 477 2144 483 2256
rect 525 2184 531 2297
rect 557 2284 563 2436
rect 573 2404 579 2436
rect 461 2124 467 2136
rect 493 2124 499 2156
rect 589 2144 595 2576
rect 605 2524 611 2676
rect 621 2544 627 2716
rect 877 2684 883 2696
rect 941 2684 947 2936
rect 957 2744 963 2936
rect 733 2464 739 2636
rect 781 2564 787 2676
rect 845 2584 851 2656
rect 925 2644 931 2676
rect 941 2624 947 2656
rect 605 2324 611 2356
rect 653 2324 659 2336
rect 621 2204 627 2236
rect 637 2183 643 2256
rect 621 2177 643 2183
rect 525 2104 531 2136
rect 573 2104 579 2116
rect 621 2084 627 2177
rect 653 2124 659 2316
rect 733 2304 739 2436
rect 781 2384 787 2556
rect 797 2544 803 2556
rect 861 2504 867 2516
rect 845 2444 851 2496
rect 893 2484 899 2516
rect 909 2503 915 2556
rect 941 2504 947 2576
rect 909 2497 924 2503
rect 941 2284 947 2496
rect 957 2444 963 2636
rect 989 2564 995 2676
rect 1005 2664 1011 2996
rect 1133 2924 1139 2956
rect 1197 2926 1203 3036
rect 1245 2864 1251 3036
rect 1261 2984 1267 3076
rect 1053 2684 1059 2716
rect 1101 2684 1107 2836
rect 1117 2704 1123 2716
rect 1092 2677 1100 2683
rect 1037 2604 1043 2636
rect 989 2544 995 2556
rect 1005 2544 1011 2556
rect 1101 2544 1107 2636
rect 973 2504 979 2516
rect 1037 2504 1043 2516
rect 1069 2484 1075 2516
rect 1101 2504 1107 2516
rect 1117 2483 1123 2696
rect 1293 2684 1299 2876
rect 1309 2723 1315 3316
rect 1325 3004 1331 3356
rect 1357 3224 1363 3236
rect 1357 3144 1363 3216
rect 1405 3144 1411 3236
rect 1485 3184 1491 3296
rect 1533 3244 1539 3318
rect 1581 3184 1587 3276
rect 1597 3224 1603 3296
rect 1613 3284 1619 3316
rect 1677 3284 1683 3316
rect 1693 3163 1699 3316
rect 1709 3183 1715 3336
rect 1725 3324 1731 3336
rect 1736 3206 1742 3214
rect 1750 3206 1756 3214
rect 1764 3206 1770 3214
rect 1778 3206 1784 3214
rect 1805 3204 1811 3636
rect 1837 3624 1843 3836
rect 1853 3784 1859 3837
rect 1885 3784 1891 3856
rect 1901 3744 1907 3756
rect 1933 3724 1939 3836
rect 1965 3764 1971 3876
rect 2093 3784 2099 3856
rect 2013 3584 2019 3756
rect 2029 3584 2035 3736
rect 2093 3724 2099 3776
rect 2205 3704 2211 3836
rect 2221 3744 2227 3756
rect 2237 3744 2243 4116
rect 2317 4064 2323 4136
rect 2269 3904 2275 3996
rect 2317 3944 2323 4056
rect 2333 4024 2339 4116
rect 2365 4104 2371 4296
rect 2413 4224 2419 4296
rect 2573 4284 2579 4796
rect 2589 4704 2595 4716
rect 2669 4704 2675 4796
rect 2733 4702 2739 4736
rect 2765 4684 2771 4696
rect 2797 4643 2803 4676
rect 2781 4637 2803 4643
rect 2589 4564 2595 4636
rect 2781 4584 2787 4637
rect 2637 4537 2675 4543
rect 2637 4524 2643 4537
rect 2669 4524 2675 4537
rect 2653 4504 2659 4516
rect 2685 4504 2691 4556
rect 2749 4524 2755 4556
rect 2797 4504 2803 4536
rect 2813 4524 2819 4596
rect 2829 4584 2835 4696
rect 2845 4684 2851 4716
rect 3117 4704 3123 4716
rect 2973 4684 2979 4696
rect 2861 4564 2867 4636
rect 3021 4603 3027 4676
rect 3021 4597 3043 4603
rect 3037 4564 3043 4597
rect 2829 4504 2835 4556
rect 3085 4544 3091 4636
rect 3149 4544 3155 4797
rect 3165 4704 3171 4796
rect 3197 4724 3203 4836
rect 3197 4704 3203 4716
rect 3165 4664 3171 4696
rect 3213 4544 3219 4876
rect 3277 4644 3283 4936
rect 3341 4904 3347 4956
rect 3373 4924 3379 5076
rect 3389 4984 3395 5080
rect 3437 4984 3443 5096
rect 3485 5064 3491 5236
rect 3549 5224 3555 5256
rect 3597 5204 3603 5296
rect 3661 5264 3667 5336
rect 3709 5304 3715 5416
rect 3869 5364 3875 5417
rect 3917 5384 3923 5476
rect 4093 5464 4099 5476
rect 4205 5464 4211 5497
rect 4269 5484 4275 5596
rect 4253 5464 4259 5476
rect 4013 5364 4019 5396
rect 3773 5326 3779 5356
rect 3517 5084 3523 5116
rect 3549 5104 3555 5116
rect 3533 5097 3548 5103
rect 3501 5064 3507 5076
rect 3389 4904 3395 4956
rect 3421 4944 3427 4956
rect 3293 4784 3299 4896
rect 3469 4864 3475 4896
rect 3533 4884 3539 5097
rect 3581 5084 3587 5096
rect 3549 4924 3555 5076
rect 3565 5004 3571 5076
rect 3661 5064 3667 5096
rect 3613 4984 3619 5056
rect 3581 4944 3587 4956
rect 3613 4944 3619 4976
rect 3549 4904 3555 4916
rect 3565 4904 3571 4916
rect 3405 4684 3411 4856
rect 3485 4704 3491 4876
rect 3549 4784 3555 4836
rect 3565 4704 3571 4896
rect 3597 4744 3603 4836
rect 3588 4717 3596 4723
rect 3549 4697 3564 4703
rect 3245 4584 3251 4616
rect 3272 4606 3278 4614
rect 3286 4606 3292 4614
rect 3300 4606 3306 4614
rect 3314 4606 3320 4614
rect 2861 4524 2867 4536
rect 3037 4504 3043 4518
rect 2669 4484 2675 4496
rect 2909 4484 2915 4496
rect 2797 4384 2803 4476
rect 2925 4384 2931 4496
rect 2429 4204 2435 4276
rect 2477 4144 2483 4236
rect 2493 4164 2499 4276
rect 2541 4184 2547 4196
rect 2589 4184 2595 4216
rect 2669 4184 2675 4316
rect 2813 4304 2819 4356
rect 2948 4317 2963 4323
rect 2957 4304 2963 4317
rect 3133 4304 3139 4476
rect 3197 4444 3203 4516
rect 3229 4484 3235 4496
rect 3261 4444 3267 4516
rect 2685 4164 2691 4256
rect 2701 4204 2707 4296
rect 2381 3984 2387 4016
rect 2413 3924 2419 3936
rect 2429 3924 2435 4036
rect 2445 3984 2451 4116
rect 2301 3884 2307 3916
rect 2429 3904 2435 3916
rect 2388 3897 2403 3903
rect 2349 3884 2355 3896
rect 2253 3784 2259 3816
rect 2317 3783 2323 3836
rect 2365 3784 2371 3876
rect 2397 3784 2403 3897
rect 2445 3864 2451 3876
rect 2301 3777 2323 3783
rect 2301 3724 2307 3777
rect 2221 3704 2227 3716
rect 2349 3704 2355 3736
rect 2381 3724 2387 3756
rect 2397 3704 2403 3756
rect 2445 3704 2451 3736
rect 2461 3724 2467 3776
rect 2477 3724 2483 4036
rect 2525 4024 2531 4156
rect 2541 3983 2547 4036
rect 2541 3977 2563 3983
rect 2525 3904 2531 3936
rect 2541 3904 2547 3956
rect 2557 3924 2563 3977
rect 2573 3964 2579 4076
rect 2509 3883 2515 3896
rect 2557 3884 2563 3916
rect 2589 3903 2595 4116
rect 2605 4024 2611 4096
rect 2580 3897 2604 3903
rect 2509 3877 2531 3883
rect 2493 3784 2499 3876
rect 2525 3784 2531 3877
rect 2589 3857 2604 3863
rect 2509 3744 2515 3756
rect 2589 3744 2595 3857
rect 2605 3724 2611 3736
rect 2317 3584 2323 3676
rect 1837 3364 1843 3376
rect 1709 3177 1731 3183
rect 1693 3157 1715 3163
rect 1341 3084 1347 3096
rect 1437 3064 1443 3136
rect 1565 3124 1571 3136
rect 1613 3084 1619 3116
rect 1501 3064 1507 3076
rect 1517 3064 1523 3076
rect 1613 3064 1619 3076
rect 1357 2944 1363 3036
rect 1405 3004 1411 3036
rect 1565 2944 1571 2996
rect 1645 2944 1651 3116
rect 1709 3084 1715 3157
rect 1725 3084 1731 3177
rect 1837 3124 1843 3356
rect 1853 3304 1859 3536
rect 1885 3502 1891 3516
rect 2157 3502 2163 3516
rect 2301 3484 2307 3516
rect 2317 3484 2323 3556
rect 2397 3484 2403 3576
rect 2477 3524 2483 3716
rect 2557 3704 2563 3716
rect 2621 3584 2627 4156
rect 2717 4124 2723 4236
rect 2781 4224 2787 4256
rect 2669 4104 2675 4116
rect 2637 3984 2643 3996
rect 2669 3884 2675 3916
rect 2685 3904 2691 3936
rect 2701 3924 2707 3956
rect 2733 3944 2739 4156
rect 2813 4144 2819 4276
rect 2829 4244 2835 4276
rect 2877 4204 2883 4236
rect 2925 4224 2931 4296
rect 2884 4177 2915 4183
rect 2909 4164 2915 4177
rect 2765 4084 2771 4096
rect 2765 4004 2771 4076
rect 2781 4064 2787 4096
rect 2692 3897 2707 3903
rect 2701 3864 2707 3897
rect 2781 3884 2787 4016
rect 2733 3784 2739 3856
rect 2749 3804 2755 3856
rect 2781 3744 2787 3876
rect 2797 3864 2803 3876
rect 2797 3744 2803 3836
rect 2781 3704 2787 3736
rect 2797 3644 2803 3736
rect 2813 3724 2819 4116
rect 2909 4104 2915 4136
rect 2845 3804 2851 3836
rect 2845 3764 2851 3796
rect 2845 3703 2851 3736
rect 2861 3724 2867 3796
rect 2877 3744 2883 4076
rect 2909 3844 2915 4096
rect 2925 3864 2931 4196
rect 3021 4184 3027 4236
rect 3053 4224 3059 4256
rect 3069 4244 3075 4276
rect 3149 4244 3155 4296
rect 3053 4164 3059 4196
rect 3117 4164 3123 4216
rect 2989 4144 2995 4156
rect 2957 3924 2963 4036
rect 2989 4004 2995 4116
rect 3053 3984 3059 4136
rect 3085 4044 3091 4096
rect 3085 3924 3091 4036
rect 3133 3984 3139 4116
rect 3165 3944 3171 4436
rect 3309 4384 3315 4496
rect 3293 4244 3299 4296
rect 3325 4264 3331 4556
rect 3405 4543 3411 4676
rect 3421 4564 3427 4596
rect 3501 4584 3507 4676
rect 3549 4664 3555 4697
rect 3405 4537 3420 4543
rect 3549 4543 3555 4656
rect 3581 4564 3587 4596
rect 3597 4584 3603 4716
rect 3629 4684 3635 4736
rect 3645 4724 3651 4996
rect 3677 4924 3683 5076
rect 3693 5004 3699 5076
rect 3709 4884 3715 5296
rect 3757 5124 3763 5136
rect 3789 5104 3795 5116
rect 3725 5084 3731 5096
rect 3741 5084 3747 5096
rect 3805 4984 3811 5156
rect 3821 4984 3827 5316
rect 3885 5104 3891 5316
rect 3917 5304 3923 5356
rect 4061 5344 4067 5396
rect 4125 5343 4131 5456
rect 4173 5424 4179 5456
rect 4116 5337 4131 5343
rect 4093 5324 4099 5336
rect 4141 5324 4147 5356
rect 4205 5344 4211 5376
rect 4157 5324 4163 5336
rect 3981 5304 3987 5316
rect 4221 5304 4227 5336
rect 4237 5324 4243 5436
rect 4269 5404 4275 5476
rect 4285 5364 4291 5476
rect 4301 5384 4307 5436
rect 4301 5363 4307 5376
rect 4301 5357 4316 5363
rect 4333 5344 4339 5416
rect 4349 5344 4355 5516
rect 4365 5504 4371 5636
rect 4381 5604 4387 5756
rect 4493 5703 4499 5736
rect 4509 5724 4515 5776
rect 4765 5757 4780 5763
rect 4525 5724 4531 5736
rect 4493 5697 4515 5703
rect 4509 5684 4515 5697
rect 4388 5597 4403 5603
rect 4397 5544 4403 5597
rect 4493 5584 4499 5676
rect 4589 5564 4595 5756
rect 4765 5643 4771 5757
rect 4756 5637 4771 5643
rect 4621 5584 4627 5636
rect 4381 5504 4387 5516
rect 4397 5484 4403 5536
rect 4413 5524 4419 5556
rect 4557 5524 4563 5556
rect 4461 5464 4467 5476
rect 3901 5204 3907 5236
rect 3901 5084 3907 5096
rect 3741 4964 3747 4976
rect 3645 4684 3651 4716
rect 3677 4684 3683 4856
rect 3741 4784 3747 4918
rect 3812 4897 3827 4903
rect 3821 4884 3827 4897
rect 3709 4704 3715 4776
rect 3805 4703 3811 4876
rect 3837 4804 3843 5056
rect 3917 5044 3923 5296
rect 3981 5244 3987 5256
rect 3869 4924 3875 5036
rect 3885 4964 3891 5036
rect 3901 4964 3907 5016
rect 3821 4724 3827 4756
rect 3805 4697 3827 4703
rect 3773 4684 3779 4696
rect 3677 4664 3683 4676
rect 3757 4664 3763 4676
rect 3693 4584 3699 4616
rect 3540 4537 3555 4543
rect 3437 4384 3443 4476
rect 3517 4384 3523 4476
rect 3453 4304 3459 4336
rect 3533 4304 3539 4336
rect 3272 4206 3278 4214
rect 3286 4206 3292 4214
rect 3300 4206 3306 4214
rect 3314 4206 3320 4214
rect 3181 4164 3187 4176
rect 3213 4144 3219 4196
rect 3389 4184 3395 4296
rect 3437 4284 3443 4296
rect 3437 4264 3443 4276
rect 3149 3902 3155 3916
rect 3197 3904 3203 4096
rect 3213 3964 3219 4036
rect 3309 3924 3315 4076
rect 3325 4024 3331 4116
rect 2957 3884 2963 3896
rect 3053 3884 3059 3896
rect 2925 3764 2931 3836
rect 2941 3784 2947 3796
rect 2973 3784 2979 3876
rect 3005 3864 3011 3876
rect 3037 3804 3043 3876
rect 3117 3864 3123 3876
rect 3053 3764 3059 3856
rect 3149 3824 3155 3856
rect 3181 3784 3187 3896
rect 3341 3884 3347 4136
rect 3485 4124 3491 4296
rect 3533 4184 3539 4276
rect 3565 4204 3571 4556
rect 3645 4484 3651 4556
rect 3725 4524 3731 4596
rect 3821 4564 3827 4697
rect 3853 4663 3859 4916
rect 3885 4784 3891 4896
rect 3869 4684 3875 4696
rect 3917 4683 3923 4836
rect 3949 4824 3955 5116
rect 3981 5104 3987 5236
rect 4013 5102 4019 5136
rect 4141 5124 4147 5236
rect 4333 5184 4339 5336
rect 4413 5323 4419 5436
rect 4493 5424 4499 5496
rect 4541 5484 4547 5516
rect 4557 5464 4563 5496
rect 4733 5484 4739 5576
rect 4621 5384 4627 5476
rect 4733 5344 4739 5476
rect 4749 5424 4755 5456
rect 4765 5363 4771 5637
rect 4808 5606 4814 5614
rect 4822 5606 4828 5614
rect 4836 5606 4842 5614
rect 4850 5606 4856 5614
rect 4973 5584 4979 5736
rect 4973 5564 4979 5576
rect 4788 5517 4803 5523
rect 4797 5484 4803 5517
rect 4989 5523 4995 5676
rect 5005 5664 5011 5716
rect 5021 5544 5027 5776
rect 5037 5764 5043 5776
rect 6141 5764 6147 5776
rect 5053 5664 5059 5756
rect 5453 5744 5459 5756
rect 4989 5517 5004 5523
rect 4829 5484 4835 5496
rect 4797 5384 4803 5476
rect 4893 5464 4899 5476
rect 4813 5364 4819 5396
rect 4925 5384 4931 5516
rect 4941 5504 4947 5516
rect 4973 5424 4979 5496
rect 4989 5484 4995 5517
rect 4749 5357 4771 5363
rect 4404 5317 4419 5323
rect 4381 5184 4387 5296
rect 4445 5184 4451 5236
rect 4205 5102 4211 5116
rect 4557 5104 4563 5316
rect 4477 5084 4483 5096
rect 3981 4984 3987 5076
rect 4141 5044 4147 5056
rect 3981 4964 3987 4976
rect 4221 4964 4227 5076
rect 4413 5044 4419 5056
rect 4157 4924 4163 4956
rect 4109 4824 4115 4836
rect 3997 4704 4003 4716
rect 3981 4684 3987 4696
rect 3917 4677 3939 4683
rect 3853 4657 3875 4663
rect 3741 4503 3747 4536
rect 3789 4504 3795 4516
rect 3741 4497 3756 4503
rect 3661 4302 3667 4436
rect 3741 4384 3747 4497
rect 3805 4304 3811 4496
rect 3821 4484 3827 4536
rect 3853 4504 3859 4536
rect 3869 4444 3875 4657
rect 3917 4644 3923 4656
rect 3917 4584 3923 4596
rect 3901 4544 3907 4576
rect 3917 4524 3923 4536
rect 3917 4504 3923 4516
rect 3837 4363 3843 4436
rect 3821 4357 3843 4363
rect 3613 4244 3619 4296
rect 3725 4244 3731 4256
rect 3757 4244 3763 4256
rect 3805 4244 3811 4276
rect 3501 4144 3507 4156
rect 3213 3784 3219 3876
rect 3341 3864 3347 3876
rect 2845 3697 2860 3703
rect 2893 3684 2899 3716
rect 1885 3264 1891 3456
rect 2013 3424 2019 3436
rect 1949 3384 1955 3396
rect 1933 3364 1939 3376
rect 1901 3324 1907 3356
rect 2141 3344 2147 3476
rect 2429 3404 2435 3476
rect 2477 3464 2483 3496
rect 2493 3464 2499 3556
rect 2589 3484 2595 3536
rect 2605 3504 2611 3556
rect 2669 3504 2675 3636
rect 2749 3464 2755 3516
rect 2765 3484 2771 3636
rect 2797 3524 2803 3576
rect 2893 3544 2899 3676
rect 2909 3504 2915 3576
rect 2925 3564 2931 3756
rect 3197 3744 3203 3756
rect 2957 3684 2963 3696
rect 2989 3584 2995 3716
rect 3213 3697 3228 3703
rect 3037 3584 3043 3636
rect 3197 3584 3203 3676
rect 2925 3504 2931 3536
rect 2941 3524 2947 3556
rect 2989 3504 2995 3536
rect 3053 3524 3059 3576
rect 3213 3524 3219 3697
rect 3245 3683 3251 3836
rect 3272 3806 3278 3814
rect 3286 3806 3292 3814
rect 3300 3806 3306 3814
rect 3314 3806 3320 3814
rect 3373 3784 3379 3916
rect 3389 3904 3395 3996
rect 3421 3824 3427 4036
rect 3469 4004 3475 4116
rect 3469 3904 3475 3996
rect 3501 3984 3507 4136
rect 3533 4104 3539 4176
rect 3533 4024 3539 4096
rect 3549 3924 3555 3976
rect 3501 3917 3539 3923
rect 3501 3904 3507 3917
rect 3533 3904 3539 3917
rect 3229 3677 3251 3683
rect 3133 3484 3139 3496
rect 2669 3444 2675 3456
rect 2765 3444 2771 3476
rect 2749 3424 2755 3436
rect 1885 3124 1891 3216
rect 1741 3104 1747 3116
rect 1693 2964 1699 3036
rect 1709 3004 1715 3076
rect 1821 3064 1827 3096
rect 1885 3084 1891 3116
rect 1981 3104 1987 3316
rect 2013 3264 2019 3336
rect 2045 3326 2051 3336
rect 2141 3284 2147 3336
rect 2253 3304 2259 3316
rect 2013 3144 2019 3236
rect 1709 2944 1715 2956
rect 1389 2744 1395 2936
rect 1581 2924 1587 2936
rect 1629 2924 1635 2936
rect 1549 2784 1555 2836
rect 1421 2724 1427 2736
rect 1309 2717 1331 2723
rect 1229 2564 1235 2676
rect 1293 2584 1299 2676
rect 1229 2544 1235 2556
rect 1309 2544 1315 2576
rect 1101 2477 1123 2483
rect 1037 2324 1043 2436
rect 1053 2324 1059 2356
rect 1069 2344 1075 2436
rect 1101 2323 1107 2477
rect 1117 2364 1123 2436
rect 1117 2324 1123 2336
rect 1101 2317 1116 2323
rect 973 2302 979 2316
rect 1133 2304 1139 2496
rect 1149 2484 1155 2536
rect 1149 2343 1155 2476
rect 1165 2384 1171 2516
rect 1181 2404 1187 2516
rect 1229 2504 1235 2536
rect 1149 2337 1171 2343
rect 749 2124 755 2196
rect 813 2164 819 2276
rect 1005 2264 1011 2276
rect 1005 2164 1011 2256
rect 1133 2184 1139 2276
rect 1149 2164 1155 2316
rect 1165 2284 1171 2337
rect 1261 2324 1267 2336
rect 1245 2317 1260 2323
rect 1181 2304 1187 2316
rect 1213 2284 1219 2316
rect 1149 2124 1155 2136
rect 669 2084 675 2096
rect 349 1924 355 1936
rect 429 1904 435 2036
rect 637 1944 643 2036
rect 685 1984 691 2116
rect 1197 2104 1203 2276
rect 1245 2264 1251 2317
rect 1245 2144 1251 2216
rect 1261 2123 1267 2236
rect 1277 2164 1283 2456
rect 1293 2164 1299 2276
rect 1325 2184 1331 2717
rect 1437 2684 1443 2736
rect 1389 2564 1395 2576
rect 1341 2544 1347 2556
rect 1405 2524 1411 2676
rect 1453 2544 1459 2756
rect 1501 2584 1507 2596
rect 1517 2564 1523 2576
rect 1469 2504 1475 2516
rect 1485 2484 1491 2556
rect 1517 2504 1523 2556
rect 1565 2544 1571 2676
rect 1613 2624 1619 2696
rect 1613 2604 1619 2616
rect 1629 2584 1635 2676
rect 1597 2544 1603 2576
rect 1613 2504 1619 2516
rect 1629 2504 1635 2536
rect 1661 2524 1667 2576
rect 1677 2544 1683 2676
rect 1693 2664 1699 2696
rect 1709 2663 1715 2936
rect 1725 2904 1731 2976
rect 1805 2944 1811 3036
rect 1837 2984 1843 3076
rect 1757 2924 1763 2936
rect 1869 2923 1875 3036
rect 1892 2937 1907 2943
rect 1901 2924 1907 2937
rect 1917 2937 1932 2943
rect 1869 2917 1884 2923
rect 1805 2884 1811 2916
rect 1853 2904 1859 2916
rect 1736 2806 1742 2814
rect 1750 2806 1756 2814
rect 1764 2806 1770 2814
rect 1778 2806 1784 2814
rect 1709 2657 1724 2663
rect 1773 2604 1779 2716
rect 1837 2684 1843 2696
rect 1773 2564 1779 2596
rect 1421 2384 1427 2436
rect 1341 2264 1347 2376
rect 1389 2304 1395 2316
rect 1437 2304 1443 2316
rect 1357 2284 1363 2296
rect 1348 2257 1363 2263
rect 1341 2184 1347 2236
rect 1277 2144 1283 2156
rect 1293 2144 1299 2156
rect 1252 2117 1267 2123
rect 909 1984 915 2076
rect 93 1864 99 1876
rect 157 1764 163 1856
rect 173 1764 179 1796
rect 45 1584 51 1716
rect 13 1344 19 1476
rect 29 1464 35 1536
rect 45 1504 51 1536
rect 77 1524 83 1736
rect 93 1584 99 1716
rect 93 1544 99 1576
rect 109 1524 115 1716
rect 173 1704 179 1716
rect 77 1484 83 1516
rect 125 1504 131 1676
rect 141 1504 147 1516
rect 157 1504 163 1676
rect 173 1524 179 1696
rect 221 1564 227 1896
rect 493 1884 499 1894
rect 461 1864 467 1876
rect 269 1824 275 1856
rect 301 1744 307 1856
rect 333 1764 339 1856
rect 429 1784 435 1856
rect 589 1784 595 1796
rect 525 1764 531 1776
rect 605 1764 611 1796
rect 621 1784 627 1836
rect 637 1804 643 1916
rect 653 1904 659 1956
rect 813 1917 828 1923
rect 765 1904 771 1916
rect 797 1904 803 1916
rect 685 1897 700 1903
rect 221 1484 227 1496
rect 77 1356 83 1456
rect 109 1344 115 1476
rect 125 1364 131 1456
rect 173 1364 179 1436
rect 125 1324 131 1356
rect 141 1324 147 1336
rect 13 964 19 1036
rect 125 984 131 1096
rect 173 1084 179 1276
rect 269 1264 275 1476
rect 285 1464 291 1556
rect 301 1324 307 1736
rect 317 1504 323 1536
rect 397 1504 403 1556
rect 333 1484 339 1496
rect 301 1284 307 1316
rect 349 1124 355 1436
rect 381 1384 387 1476
rect 397 1364 403 1496
rect 413 1484 419 1516
rect 445 1504 451 1696
rect 461 1544 467 1636
rect 429 1384 435 1496
rect 477 1444 483 1716
rect 541 1684 547 1756
rect 548 1497 563 1503
rect 493 1484 499 1496
rect 525 1484 531 1496
rect 557 1464 563 1497
rect 381 1324 387 1356
rect 429 1324 435 1376
rect 381 1304 387 1316
rect 445 1304 451 1356
rect 461 1344 467 1356
rect 493 1324 499 1436
rect 525 1384 531 1456
rect 557 1384 563 1436
rect 365 1284 371 1296
rect 365 1184 371 1256
rect 365 1103 371 1156
rect 461 1124 467 1316
rect 493 1264 499 1296
rect 429 1104 435 1116
rect 356 1097 371 1103
rect 205 1044 211 1076
rect 13 884 19 956
rect 45 944 51 956
rect 109 944 115 976
rect 141 944 147 956
rect 157 924 163 936
rect 29 844 35 916
rect 173 904 179 916
rect 77 864 83 896
rect 29 744 35 836
rect 29 704 35 736
rect 13 684 19 696
rect 61 604 67 716
rect 77 704 83 856
rect 125 684 131 756
rect 141 724 147 876
rect 221 724 227 1036
rect 237 984 243 1036
rect 301 964 307 1076
rect 237 784 243 956
rect 317 943 323 1036
rect 413 1004 419 1076
rect 308 937 323 943
rect 269 784 275 916
rect 253 724 259 736
rect 13 584 19 596
rect 93 524 99 676
rect 141 544 147 716
rect 221 684 227 716
rect 301 704 307 916
rect 317 884 323 896
rect 365 864 371 916
rect 445 903 451 916
rect 436 897 451 903
rect 372 857 387 863
rect 301 584 307 696
rect 173 544 179 576
rect 285 544 291 556
rect 173 284 179 536
rect 333 504 339 556
rect 349 524 355 636
rect 365 564 371 776
rect 381 684 387 857
rect 397 704 403 776
rect 413 743 419 836
rect 413 737 435 743
rect 429 704 435 737
rect 461 724 467 1036
rect 509 964 515 1016
rect 541 964 547 1376
rect 573 1344 579 1456
rect 605 1364 611 1676
rect 621 1504 627 1776
rect 637 1744 643 1756
rect 669 1744 675 1896
rect 685 1704 691 1897
rect 813 1884 819 1917
rect 845 1904 851 1916
rect 797 1877 812 1883
rect 701 1783 707 1876
rect 701 1777 716 1783
rect 717 1744 723 1776
rect 701 1484 707 1736
rect 765 1724 771 1736
rect 781 1724 787 1756
rect 797 1744 803 1877
rect 861 1844 867 1936
rect 909 1864 915 1896
rect 829 1750 835 1776
rect 893 1744 899 1816
rect 909 1764 915 1836
rect 941 1824 947 1856
rect 957 1764 963 1876
rect 941 1757 956 1763
rect 893 1724 899 1736
rect 733 1504 739 1636
rect 909 1504 915 1596
rect 557 1304 563 1336
rect 573 1284 579 1316
rect 573 1104 579 1276
rect 605 1183 611 1356
rect 637 1344 643 1476
rect 589 1177 611 1183
rect 557 1083 563 1096
rect 557 1077 579 1083
rect 573 984 579 1077
rect 589 1024 595 1177
rect 557 964 563 976
rect 381 524 387 596
rect 397 584 403 676
rect 509 644 515 956
rect 589 904 595 936
rect 525 764 531 836
rect 605 784 611 996
rect 621 864 627 1296
rect 653 1084 659 1436
rect 669 1364 675 1396
rect 685 1384 691 1476
rect 893 1404 899 1436
rect 669 1124 675 1316
rect 749 1184 755 1316
rect 861 1204 867 1236
rect 909 1164 915 1496
rect 925 1404 931 1756
rect 941 1744 947 1757
rect 973 1744 979 1896
rect 989 1844 995 1916
rect 1005 1904 1011 1916
rect 1069 1904 1075 2076
rect 1293 2064 1299 2136
rect 1309 2124 1315 2136
rect 1309 1984 1315 2116
rect 1085 1904 1091 1916
rect 1165 1904 1171 1916
rect 1037 1784 1043 1876
rect 1053 1744 1059 1756
rect 1069 1744 1075 1876
rect 1117 1864 1123 1896
rect 941 1584 947 1736
rect 957 1704 963 1736
rect 1005 1704 1011 1716
rect 973 1484 979 1496
rect 1005 1363 1011 1696
rect 1053 1684 1059 1736
rect 1085 1724 1091 1836
rect 1133 1784 1139 1896
rect 1181 1884 1187 1896
rect 1197 1884 1203 1896
rect 1229 1744 1235 1976
rect 1325 1924 1331 2176
rect 1357 2144 1363 2257
rect 1373 2184 1379 2296
rect 1469 2284 1475 2336
rect 1405 2244 1411 2276
rect 1389 2084 1395 2136
rect 1421 2103 1427 2196
rect 1437 2104 1443 2276
rect 1485 2184 1491 2396
rect 1517 2344 1523 2476
rect 1565 2364 1571 2436
rect 1549 2323 1555 2356
rect 1549 2317 1571 2323
rect 1565 2304 1571 2317
rect 1645 2264 1651 2276
rect 1501 2164 1507 2236
rect 1613 2164 1619 2256
rect 1677 2204 1683 2536
rect 1741 2524 1747 2536
rect 1693 2484 1699 2496
rect 1789 2484 1795 2556
rect 1821 2484 1827 2616
rect 1837 2524 1843 2536
rect 1853 2524 1859 2776
rect 1869 2624 1875 2716
rect 1885 2544 1891 2736
rect 1917 2704 1923 2937
rect 1949 2884 1955 2916
rect 1949 2704 1955 2876
rect 1949 2684 1955 2696
rect 1997 2664 2003 3116
rect 2013 3084 2019 3096
rect 2013 2984 2019 3076
rect 2013 2924 2019 2976
rect 2029 2944 2035 3076
rect 2045 2924 2051 2956
rect 2077 2744 2083 3116
rect 2109 3084 2115 3236
rect 2141 3084 2147 3276
rect 2173 3084 2179 3236
rect 2189 3104 2195 3116
rect 2317 3064 2323 3076
rect 2173 2944 2179 3056
rect 2365 2984 2371 3096
rect 2381 2984 2387 3316
rect 2445 3284 2451 3336
rect 2461 3284 2467 3316
rect 2477 3304 2483 3376
rect 2509 3303 2515 3356
rect 2589 3344 2595 3356
rect 2541 3304 2547 3316
rect 2500 3297 2515 3303
rect 2413 3164 2419 3236
rect 2493 3184 2499 3276
rect 2541 3184 2547 3296
rect 2557 3164 2563 3336
rect 2477 3124 2483 3156
rect 2509 3124 2515 3136
rect 2445 3104 2451 3116
rect 2333 2924 2339 2976
rect 2413 2940 2419 3076
rect 2493 2984 2499 3096
rect 2557 3064 2563 3156
rect 2573 3104 2579 3316
rect 2589 3064 2595 3076
rect 2605 3044 2611 3336
rect 2621 3244 2627 3356
rect 2701 3344 2707 3356
rect 2749 3304 2755 3376
rect 2765 3364 2771 3436
rect 2797 3384 2803 3436
rect 2628 3237 2643 3243
rect 2637 3104 2643 3237
rect 2653 3104 2659 3116
rect 2445 2944 2451 2976
rect 2461 2924 2467 2976
rect 2573 2944 2579 2976
rect 2589 2944 2595 3036
rect 2605 2964 2611 3036
rect 2621 2944 2627 2956
rect 2637 2943 2643 3096
rect 2628 2937 2643 2943
rect 2653 2904 2659 3036
rect 2045 2704 2051 2716
rect 2061 2684 2067 2696
rect 1933 2544 1939 2556
rect 1949 2524 1955 2656
rect 1965 2584 1971 2636
rect 1997 2564 2003 2596
rect 2029 2584 2035 2656
rect 2061 2564 2067 2656
rect 2077 2624 2083 2696
rect 1853 2504 1859 2516
rect 1901 2484 1907 2516
rect 1917 2504 1923 2516
rect 1837 2464 1843 2476
rect 1885 2464 1891 2476
rect 1736 2406 1742 2414
rect 1750 2406 1756 2414
rect 1764 2406 1770 2414
rect 1778 2406 1784 2414
rect 1901 2324 1907 2436
rect 2029 2304 2035 2356
rect 2061 2324 2067 2376
rect 2093 2264 2099 2696
rect 2109 2504 2115 2736
rect 2141 2684 2147 2776
rect 2125 2544 2131 2616
rect 2253 2604 2259 2636
rect 2109 2383 2115 2496
rect 2109 2377 2124 2383
rect 2109 2264 2115 2276
rect 1581 2144 1587 2156
rect 1661 2124 1667 2156
rect 1789 2144 1795 2156
rect 1412 2097 1427 2103
rect 1245 1904 1251 1916
rect 1341 1904 1347 2036
rect 1309 1784 1315 1836
rect 1117 1704 1123 1716
rect 1165 1584 1171 1676
rect 1021 1504 1027 1516
rect 1069 1504 1075 1576
rect 1053 1384 1059 1496
rect 1101 1403 1107 1556
rect 1197 1504 1203 1516
rect 1229 1464 1235 1476
rect 1085 1397 1107 1403
rect 1085 1364 1091 1397
rect 1101 1364 1107 1376
rect 1005 1357 1020 1363
rect 1021 1344 1027 1356
rect 1149 1344 1155 1396
rect 1165 1364 1171 1456
rect 1261 1384 1267 1496
rect 1277 1344 1283 1436
rect 1293 1384 1299 1476
rect 1309 1444 1315 1456
rect 1325 1423 1331 1656
rect 1341 1564 1347 1896
rect 1357 1884 1363 1996
rect 1405 1904 1411 1956
rect 1421 1884 1427 2097
rect 1357 1504 1363 1856
rect 1421 1844 1427 1876
rect 1373 1744 1379 1756
rect 1421 1744 1427 1836
rect 1453 1764 1459 1956
rect 1469 1904 1475 1916
rect 1485 1844 1491 1856
rect 1389 1684 1395 1696
rect 1453 1584 1459 1696
rect 1501 1664 1507 2116
rect 1533 1724 1539 1736
rect 1469 1504 1475 1516
rect 1357 1484 1363 1496
rect 1389 1477 1404 1483
rect 1341 1464 1347 1476
rect 1389 1444 1395 1477
rect 1309 1417 1331 1423
rect 1309 1384 1315 1417
rect 1341 1364 1347 1396
rect 1325 1344 1331 1356
rect 1341 1344 1347 1356
rect 1421 1344 1427 1456
rect 637 1057 652 1063
rect 637 964 643 1057
rect 653 1044 659 1056
rect 701 1044 707 1096
rect 717 1084 723 1096
rect 749 1084 755 1096
rect 941 1084 947 1096
rect 669 984 675 1036
rect 749 944 755 1016
rect 765 904 771 1016
rect 781 984 787 1076
rect 829 944 835 1016
rect 845 944 851 1076
rect 877 924 883 1076
rect 957 1024 963 1076
rect 973 1044 979 1096
rect 941 924 947 956
rect 973 943 979 1036
rect 989 1024 995 1056
rect 1005 983 1011 1336
rect 1133 1324 1139 1336
rect 1277 1304 1283 1336
rect 1437 1324 1443 1496
rect 1485 1464 1491 1476
rect 1485 1404 1491 1456
rect 1501 1444 1507 1636
rect 1549 1604 1555 2076
rect 1597 1964 1603 2036
rect 1597 1904 1603 1936
rect 1677 1884 1683 2116
rect 1805 2104 1811 2116
rect 1736 2006 1742 2014
rect 1750 2006 1756 2014
rect 1764 2006 1770 2014
rect 1778 2006 1784 2014
rect 1805 1903 1811 2096
rect 1821 2044 1827 2256
rect 1853 2164 1859 2236
rect 1869 2084 1875 2256
rect 1901 2244 1907 2256
rect 1981 2164 1987 2256
rect 2061 2124 2067 2236
rect 1885 2104 1891 2116
rect 1949 2084 1955 2096
rect 1869 1904 1875 2076
rect 1796 1897 1811 1903
rect 1597 1764 1603 1876
rect 1677 1864 1683 1876
rect 1693 1764 1699 1836
rect 1821 1744 1827 1836
rect 1837 1804 1843 1836
rect 1869 1784 1875 1896
rect 1933 1884 1939 2036
rect 1981 1904 1987 2076
rect 2141 1963 2147 2576
rect 2221 2544 2227 2556
rect 2285 2544 2291 2836
rect 2301 2784 2307 2836
rect 2365 2704 2371 2716
rect 2189 2304 2195 2436
rect 2237 2304 2243 2316
rect 2253 2304 2259 2516
rect 2173 2144 2179 2156
rect 2189 2144 2195 2296
rect 2269 2124 2275 2216
rect 2125 1957 2147 1963
rect 2125 1904 2131 1957
rect 2157 1923 2163 2116
rect 2141 1917 2163 1923
rect 1933 1744 1939 1856
rect 1693 1724 1699 1736
rect 1597 1684 1603 1718
rect 1645 1584 1651 1676
rect 1677 1624 1683 1636
rect 1736 1606 1742 1614
rect 1750 1606 1756 1614
rect 1764 1606 1770 1614
rect 1778 1606 1784 1614
rect 1581 1524 1587 1536
rect 1613 1517 1628 1523
rect 1581 1464 1587 1516
rect 1597 1464 1603 1476
rect 1469 1324 1475 1376
rect 1501 1344 1507 1436
rect 1533 1384 1539 1436
rect 1565 1323 1571 1436
rect 1597 1344 1603 1456
rect 1613 1384 1619 1517
rect 1677 1484 1683 1516
rect 1693 1504 1699 1556
rect 1709 1524 1715 1556
rect 1805 1524 1811 1716
rect 1837 1524 1843 1576
rect 1869 1563 1875 1736
rect 1853 1557 1875 1563
rect 1709 1484 1715 1496
rect 1613 1324 1619 1336
rect 1629 1324 1635 1436
rect 1645 1344 1651 1456
rect 1693 1384 1699 1476
rect 1565 1317 1580 1323
rect 1021 1144 1027 1196
rect 1021 1064 1027 1136
rect 964 937 979 943
rect 989 977 1011 983
rect 685 884 691 896
rect 861 884 867 896
rect 973 884 979 916
rect 685 702 691 716
rect 477 564 483 636
rect 429 544 435 556
rect 445 524 451 536
rect 413 504 419 516
rect 221 283 227 336
rect 237 304 243 336
rect 333 324 339 496
rect 573 444 579 556
rect 701 524 707 676
rect 813 644 819 656
rect 637 504 643 518
rect 349 344 355 356
rect 205 277 227 283
rect 20 237 35 243
rect 13 144 19 216
rect 29 164 35 237
rect 93 184 99 256
rect 205 184 211 277
rect 29 124 35 156
rect 61 124 67 136
rect 77 124 83 156
rect 141 124 147 156
rect 253 144 259 276
rect 269 264 275 276
rect 285 184 291 296
rect 333 143 339 316
rect 349 164 355 296
rect 324 137 339 143
rect 349 124 355 156
rect 237 104 243 116
rect 365 103 371 336
rect 461 304 467 436
rect 397 264 403 276
rect 429 224 435 256
rect 397 184 403 196
rect 413 104 419 136
rect 445 124 451 296
rect 509 284 515 316
rect 573 304 579 336
rect 493 277 508 283
rect 477 164 483 276
rect 477 124 483 156
rect 493 144 499 277
rect 557 184 563 276
rect 621 264 627 276
rect 589 144 595 176
rect 605 124 611 236
rect 717 184 723 216
rect 717 144 723 156
rect 653 137 668 143
rect 621 124 627 136
rect 653 124 659 137
rect 749 104 755 136
rect 765 124 771 336
rect 781 304 787 516
rect 813 504 819 636
rect 845 524 851 676
rect 989 604 995 977
rect 1021 964 1027 1056
rect 1037 944 1043 1056
rect 1069 944 1075 1236
rect 1101 1064 1107 1136
rect 1005 884 1011 896
rect 1005 784 1011 876
rect 1037 704 1043 916
rect 1085 904 1091 1056
rect 1117 1043 1123 1096
rect 1197 1064 1203 1076
rect 1101 1037 1123 1043
rect 1101 904 1107 1037
rect 1117 944 1123 1016
rect 1117 704 1123 916
rect 1133 904 1139 1036
rect 1213 964 1219 1076
rect 1229 1044 1235 1296
rect 1277 1184 1283 1276
rect 1181 904 1187 936
rect 1213 924 1219 956
rect 1245 944 1251 1116
rect 1277 1084 1283 1136
rect 1533 1123 1539 1276
rect 1581 1164 1587 1236
rect 1661 1184 1667 1296
rect 1709 1124 1715 1416
rect 1736 1206 1742 1214
rect 1750 1206 1756 1214
rect 1764 1206 1770 1214
rect 1778 1206 1784 1214
rect 1821 1184 1827 1476
rect 1853 1364 1859 1557
rect 1869 1484 1875 1536
rect 1917 1484 1923 1536
rect 2013 1484 2019 1636
rect 1948 1464 1956 1470
rect 2029 1463 2035 1716
rect 2045 1504 2051 1876
rect 2125 1844 2131 1856
rect 2045 1464 2051 1496
rect 2061 1484 2067 1796
rect 2077 1724 2083 1836
rect 2093 1684 2099 1716
rect 2013 1457 2035 1463
rect 1965 1344 1971 1376
rect 1917 1324 1923 1336
rect 1981 1304 1987 1336
rect 1533 1117 1548 1123
rect 1357 1084 1363 1096
rect 1437 1084 1443 1116
rect 1341 1064 1347 1076
rect 1389 1044 1395 1056
rect 1405 1044 1411 1076
rect 1453 1064 1459 1096
rect 1709 1084 1715 1116
rect 1757 1084 1763 1116
rect 1933 1104 1939 1156
rect 1453 1044 1459 1056
rect 1485 1044 1491 1076
rect 1293 1024 1299 1036
rect 1261 924 1267 976
rect 1293 924 1299 936
rect 1309 924 1315 996
rect 1389 944 1395 1036
rect 1405 944 1411 1036
rect 1421 1004 1427 1036
rect 1469 1004 1475 1036
rect 1485 1024 1491 1036
rect 1485 984 1491 1016
rect 1533 1004 1539 1036
rect 1597 983 1603 1036
rect 1581 977 1603 983
rect 1341 924 1347 936
rect 1229 904 1235 916
rect 1213 784 1219 896
rect 1229 744 1235 856
rect 1341 784 1347 896
rect 1293 684 1299 736
rect 1341 724 1347 776
rect 1373 744 1379 916
rect 1421 904 1427 936
rect 1421 683 1427 896
rect 1453 884 1459 956
rect 1485 944 1491 976
rect 1501 924 1507 956
rect 1549 904 1555 956
rect 1581 944 1587 977
rect 1597 924 1603 956
rect 1629 923 1635 936
rect 1613 917 1635 923
rect 1565 903 1571 916
rect 1613 903 1619 917
rect 1565 897 1619 903
rect 1645 884 1651 896
rect 1437 704 1443 836
rect 1501 764 1507 836
rect 1533 724 1539 876
rect 1581 724 1587 756
rect 1421 677 1436 683
rect 925 544 931 596
rect 1037 584 1043 676
rect 1117 564 1123 676
rect 1197 644 1203 676
rect 1229 664 1235 676
rect 1501 664 1507 676
rect 1293 644 1299 656
rect 1485 644 1491 656
rect 1245 603 1251 636
rect 1229 597 1251 603
rect 813 164 819 436
rect 861 224 867 316
rect 813 144 819 156
rect 845 144 851 176
rect 797 104 803 116
rect 877 104 883 236
rect 893 204 899 296
rect 1037 284 1043 436
rect 1133 384 1139 536
rect 1149 524 1155 556
rect 1229 483 1235 597
rect 1261 564 1267 636
rect 1325 564 1331 596
rect 1389 564 1395 636
rect 1533 583 1539 716
rect 1645 704 1651 716
rect 1661 704 1667 916
rect 1677 904 1683 1076
rect 1709 944 1715 976
rect 1725 904 1731 916
rect 1741 844 1747 1036
rect 1805 983 1811 1076
rect 1805 977 1820 983
rect 1805 964 1811 977
rect 1677 724 1683 836
rect 1709 704 1715 836
rect 1736 806 1742 814
rect 1750 806 1756 814
rect 1764 806 1770 814
rect 1778 806 1784 814
rect 1773 704 1779 716
rect 1805 704 1811 716
rect 1693 664 1699 676
rect 1581 584 1587 636
rect 1597 624 1603 656
rect 1837 644 1843 1056
rect 1981 944 1987 1076
rect 2013 1064 2019 1457
rect 2029 1384 2035 1436
rect 2061 1364 2067 1396
rect 2109 1363 2115 1436
rect 2125 1424 2131 1436
rect 2141 1384 2147 1917
rect 2173 1903 2179 2116
rect 2221 1924 2227 1936
rect 2269 1924 2275 1956
rect 2164 1897 2179 1903
rect 2173 1504 2179 1897
rect 2189 1784 2195 1856
rect 2237 1824 2243 1896
rect 2269 1764 2275 1836
rect 2205 1684 2211 1736
rect 2285 1524 2291 2436
rect 2317 2404 2323 2636
rect 2381 2584 2387 2656
rect 2365 2524 2371 2536
rect 2317 2224 2323 2256
rect 2301 2024 2307 2036
rect 2333 1964 2339 2236
rect 2349 2184 2355 2236
rect 2365 2224 2371 2496
rect 2413 2284 2419 2676
rect 2461 2564 2467 2796
rect 2669 2784 2675 3276
rect 2781 3244 2787 3356
rect 2797 3304 2803 3336
rect 2813 3244 2819 3456
rect 2877 3424 2883 3456
rect 2829 3364 2835 3396
rect 2845 3304 2851 3416
rect 2941 3384 2947 3396
rect 3005 3384 3011 3456
rect 2877 3324 2883 3376
rect 2925 3344 2931 3356
rect 2685 3084 2691 3156
rect 2717 3123 2723 3236
rect 2717 3117 2739 3123
rect 2733 3064 2739 3117
rect 2765 3084 2771 3116
rect 2797 3084 2803 3156
rect 2701 2944 2707 3056
rect 2893 3044 2899 3076
rect 2909 3064 2915 3196
rect 2941 3184 2947 3196
rect 2749 3003 2755 3036
rect 2749 2997 2771 3003
rect 2701 2904 2707 2936
rect 2765 2926 2771 2997
rect 2797 2704 2803 2936
rect 2941 2924 2947 2936
rect 2893 2884 2899 2896
rect 2909 2884 2915 2896
rect 2861 2784 2867 2796
rect 2877 2784 2883 2836
rect 2909 2704 2915 2856
rect 2957 2784 2963 3336
rect 3021 3064 3027 3476
rect 3117 3344 3123 3456
rect 3229 3340 3235 3677
rect 3277 3644 3283 3716
rect 3341 3704 3347 3716
rect 3373 3684 3379 3776
rect 3405 3704 3411 3736
rect 3437 3724 3443 3756
rect 3453 3744 3459 3856
rect 3469 3764 3475 3896
rect 3485 3764 3491 3896
rect 3517 3884 3523 3896
rect 3581 3884 3587 3896
rect 3565 3864 3571 3876
rect 3581 3844 3587 3876
rect 3501 3664 3507 3756
rect 3533 3744 3539 3816
rect 3549 3803 3555 3836
rect 3549 3797 3571 3803
rect 3565 3783 3571 3797
rect 3565 3777 3587 3783
rect 3549 3724 3555 3776
rect 3565 3744 3571 3756
rect 3581 3724 3587 3777
rect 3597 3744 3603 3856
rect 3613 3764 3619 4236
rect 3757 4164 3763 4176
rect 3709 4144 3715 4156
rect 3773 4124 3779 4156
rect 3821 4143 3827 4357
rect 3837 4324 3843 4336
rect 3869 4244 3875 4436
rect 3885 4284 3891 4336
rect 3917 4164 3923 4276
rect 3933 4144 3939 4677
rect 3949 4624 3955 4656
rect 3949 4544 3955 4576
rect 3997 4524 4003 4696
rect 4109 4684 4115 4736
rect 3949 4484 3955 4516
rect 3981 4504 3987 4516
rect 3965 4464 3971 4496
rect 3997 4484 4003 4516
rect 4013 4464 4019 4676
rect 4045 4584 4051 4670
rect 4125 4663 4131 4676
rect 4109 4657 4131 4663
rect 3972 4457 3987 4463
rect 3965 4304 3971 4436
rect 3981 4284 3987 4457
rect 4045 4404 4051 4436
rect 4013 4324 4019 4336
rect 3812 4137 3827 4143
rect 3949 4124 3955 4236
rect 3997 4144 4003 4316
rect 3693 4064 3699 4116
rect 3661 4004 3667 4036
rect 3693 3937 3811 3943
rect 3693 3924 3699 3937
rect 3645 3897 3660 3903
rect 3629 3864 3635 3876
rect 3645 3784 3651 3897
rect 3709 3844 3715 3896
rect 3741 3863 3747 3896
rect 3725 3857 3747 3863
rect 3725 3784 3731 3857
rect 3757 3764 3763 3916
rect 3773 3904 3779 3916
rect 3789 3904 3795 3916
rect 3805 3884 3811 3937
rect 3821 3924 3827 4036
rect 3844 3957 3891 3963
rect 3869 3903 3875 3936
rect 3885 3904 3891 3957
rect 3860 3897 3875 3903
rect 3789 3764 3795 3856
rect 3837 3844 3843 3876
rect 3901 3844 3907 4116
rect 3933 3904 3939 4016
rect 3629 3724 3635 3756
rect 3645 3704 3651 3716
rect 3661 3704 3667 3756
rect 3709 3744 3715 3756
rect 3709 3724 3715 3736
rect 3789 3726 3795 3736
rect 3917 3684 3923 3716
rect 3357 3544 3363 3636
rect 3437 3564 3443 3636
rect 3453 3584 3459 3636
rect 3581 3624 3587 3636
rect 3245 3504 3251 3536
rect 3357 3504 3363 3516
rect 3517 3504 3523 3576
rect 3261 3464 3267 3476
rect 3357 3464 3363 3496
rect 3389 3464 3395 3476
rect 3272 3406 3278 3414
rect 3286 3406 3292 3414
rect 3300 3406 3306 3414
rect 3314 3406 3320 3414
rect 3389 3384 3395 3456
rect 3437 3424 3443 3496
rect 3069 3084 3075 3316
rect 3117 3304 3123 3316
rect 3165 3304 3171 3336
rect 3197 3324 3203 3336
rect 3245 3143 3251 3316
rect 3341 3224 3347 3336
rect 3373 3324 3379 3356
rect 3469 3324 3475 3436
rect 3485 3324 3491 3476
rect 3501 3444 3507 3496
rect 3517 3484 3523 3496
rect 3565 3444 3571 3476
rect 3245 3137 3267 3143
rect 2989 2964 2995 2976
rect 3149 2964 3155 3096
rect 3181 2984 3187 3096
rect 3197 3084 3203 3116
rect 3261 3043 3267 3137
rect 3325 3104 3331 3136
rect 3357 3104 3363 3296
rect 3373 3284 3379 3316
rect 3501 3304 3507 3356
rect 3533 3344 3539 3436
rect 3565 3326 3571 3376
rect 3421 3124 3427 3136
rect 3469 3123 3475 3136
rect 3437 3117 3475 3123
rect 3437 3103 3443 3117
rect 3533 3104 3539 3156
rect 3613 3144 3619 3676
rect 3933 3663 3939 3696
rect 3917 3657 3939 3663
rect 3645 3424 3651 3496
rect 3661 3464 3667 3516
rect 3677 3464 3683 3476
rect 3693 3424 3699 3496
rect 3629 3304 3635 3316
rect 3661 3303 3667 3336
rect 3725 3323 3731 3536
rect 3741 3504 3747 3556
rect 3773 3524 3779 3556
rect 3853 3544 3859 3556
rect 3741 3444 3747 3456
rect 3805 3444 3811 3496
rect 3821 3484 3827 3516
rect 3853 3497 3868 3503
rect 3853 3484 3859 3497
rect 3757 3344 3763 3436
rect 3789 3344 3795 3376
rect 3821 3364 3827 3476
rect 3869 3384 3875 3416
rect 3901 3344 3907 3436
rect 3917 3384 3923 3657
rect 3965 3604 3971 4116
rect 3997 4104 4003 4136
rect 4013 4124 4019 4196
rect 4029 4184 4035 4276
rect 4045 4184 4051 4376
rect 4061 4344 4067 4636
rect 4109 4564 4115 4657
rect 4077 4444 4083 4476
rect 4109 4464 4115 4556
rect 4077 4423 4083 4436
rect 4077 4417 4099 4423
rect 4077 4324 4083 4396
rect 4093 4384 4099 4417
rect 4125 4224 4131 4516
rect 4141 4444 4147 4876
rect 4285 4704 4291 4776
rect 4157 4543 4163 4636
rect 4237 4584 4243 4596
rect 4221 4564 4227 4576
rect 4285 4544 4291 4696
rect 4333 4584 4339 5036
rect 4445 4964 4451 5056
rect 4420 4917 4435 4923
rect 4349 4804 4355 4836
rect 4349 4704 4355 4736
rect 4397 4704 4403 4836
rect 4429 4784 4435 4917
rect 4445 4764 4451 4956
rect 4605 4924 4611 5256
rect 4733 5124 4739 5136
rect 4749 5124 4755 5357
rect 4925 5344 4931 5376
rect 4989 5364 4995 5476
rect 5021 5424 5027 5496
rect 4989 5344 4995 5356
rect 4701 5084 4707 5096
rect 4660 5057 4675 5063
rect 4637 4984 4643 5036
rect 4669 4940 4675 5057
rect 4701 4984 4707 5056
rect 4749 4944 4755 4996
rect 4765 4944 4771 5336
rect 4781 5244 4787 5316
rect 4808 5206 4814 5214
rect 4822 5206 4828 5214
rect 4836 5206 4842 5214
rect 4850 5206 4856 5214
rect 4829 5144 4835 5176
rect 4877 5164 4883 5276
rect 4797 5084 4803 5116
rect 4877 5104 4883 5156
rect 4893 5144 4899 5316
rect 4909 5304 4915 5316
rect 4941 5264 4947 5316
rect 4909 5084 4915 5176
rect 5005 5124 5011 5356
rect 5053 5304 5059 5536
rect 5085 5464 5091 5736
rect 5133 5724 5139 5736
rect 5181 5704 5187 5716
rect 5213 5704 5219 5736
rect 5245 5726 5251 5736
rect 5117 5684 5123 5696
rect 5373 5684 5379 5696
rect 5389 5684 5395 5736
rect 5501 5724 5507 5736
rect 5069 5324 5075 5416
rect 5101 5384 5107 5496
rect 5133 5484 5139 5516
rect 5341 5504 5347 5676
rect 5389 5584 5395 5676
rect 5421 5644 5427 5696
rect 5469 5584 5475 5656
rect 5533 5584 5539 5636
rect 5117 5464 5123 5476
rect 5197 5424 5203 5436
rect 5117 5344 5123 5376
rect 5149 5324 5155 5416
rect 5181 5324 5187 5356
rect 4925 5104 4931 5116
rect 5085 5103 5091 5236
rect 5149 5184 5155 5236
rect 5213 5104 5219 5356
rect 5229 5344 5235 5456
rect 5245 5344 5251 5436
rect 5261 5423 5267 5496
rect 5277 5444 5283 5456
rect 5261 5417 5283 5423
rect 5229 5324 5235 5336
rect 5245 5304 5251 5336
rect 5277 5324 5283 5417
rect 5341 5364 5347 5496
rect 5437 5464 5443 5476
rect 5469 5443 5475 5496
rect 5517 5484 5523 5516
rect 5549 5484 5555 5756
rect 5565 5664 5571 5736
rect 5581 5584 5587 5756
rect 5629 5504 5635 5596
rect 5677 5484 5683 5756
rect 5709 5684 5715 5736
rect 5741 5683 5747 5756
rect 5885 5744 5891 5756
rect 5773 5684 5779 5716
rect 5789 5704 5795 5716
rect 5821 5704 5827 5716
rect 5725 5677 5747 5683
rect 5725 5624 5731 5677
rect 5741 5604 5747 5636
rect 5757 5604 5763 5656
rect 5805 5644 5811 5696
rect 5837 5664 5843 5736
rect 5853 5704 5859 5736
rect 5869 5684 5875 5716
rect 5917 5684 5923 5736
rect 5757 5504 5763 5596
rect 5789 5504 5795 5636
rect 5805 5524 5811 5556
rect 5885 5484 5891 5636
rect 5917 5604 5923 5676
rect 5508 5457 5523 5463
rect 5453 5437 5475 5443
rect 5453 5384 5459 5437
rect 5517 5364 5523 5457
rect 5549 5444 5555 5476
rect 5581 5464 5587 5476
rect 5885 5464 5891 5476
rect 5933 5444 5939 5716
rect 5949 5644 5955 5736
rect 5997 5584 6003 5616
rect 6045 5484 6051 5736
rect 6093 5724 6099 5736
rect 6157 5724 6163 5796
rect 6573 5744 6579 5756
rect 6781 5744 6787 5756
rect 7053 5744 7059 5756
rect 7165 5744 7171 5756
rect 7325 5744 7331 5756
rect 6653 5724 6659 5736
rect 6061 5664 6067 5696
rect 6093 5584 6099 5676
rect 6189 5504 6195 5576
rect 6205 5544 6211 5636
rect 6509 5504 6515 5536
rect 6589 5524 6595 5636
rect 6749 5584 6755 5716
rect 6893 5544 6899 5636
rect 6621 5504 6627 5516
rect 5949 5444 5955 5456
rect 5709 5384 5715 5436
rect 5293 5344 5299 5356
rect 5549 5344 5555 5356
rect 5277 5184 5283 5316
rect 5293 5184 5299 5336
rect 5437 5324 5443 5336
rect 5341 5284 5347 5316
rect 5421 5104 5427 5316
rect 5076 5097 5091 5103
rect 5501 5084 5507 5336
rect 5837 5326 5843 5436
rect 6125 5424 6131 5456
rect 6189 5424 6195 5456
rect 5901 5364 5907 5416
rect 5965 5364 5971 5396
rect 4781 5044 4787 5076
rect 4941 5064 4947 5076
rect 5101 5064 5107 5076
rect 4781 4984 4787 5036
rect 4605 4844 4611 4916
rect 4477 4784 4483 4836
rect 4349 4644 4355 4696
rect 4445 4644 4451 4716
rect 4477 4704 4483 4756
rect 4493 4704 4499 4776
rect 4525 4664 4531 4676
rect 4573 4664 4579 4676
rect 4589 4664 4595 4696
rect 4605 4684 4611 4696
rect 4621 4684 4627 4896
rect 4637 4744 4643 4796
rect 4733 4704 4739 4716
rect 4749 4704 4755 4876
rect 4808 4806 4814 4814
rect 4822 4806 4828 4814
rect 4836 4806 4842 4814
rect 4850 4806 4856 4814
rect 4909 4764 4915 4976
rect 5133 4964 5139 5076
rect 5517 5063 5523 5076
rect 5533 5064 5539 5116
rect 5661 5104 5667 5316
rect 5501 5057 5523 5063
rect 5229 4984 5235 5056
rect 4941 4824 4947 4918
rect 5133 4884 5139 4918
rect 5149 4784 5155 4816
rect 4829 4704 4835 4716
rect 4669 4664 4675 4696
rect 4701 4664 4707 4696
rect 4509 4644 4515 4656
rect 4157 4537 4172 4543
rect 4173 4504 4179 4516
rect 4189 4504 4195 4516
rect 4221 4364 4227 4496
rect 4253 4284 4259 4536
rect 4381 4526 4387 4596
rect 4301 4384 4307 4416
rect 4349 4384 4355 4516
rect 4317 4284 4323 4296
rect 3981 4024 3987 4096
rect 4029 3984 4035 4096
rect 4077 4064 4083 4136
rect 4061 4004 4067 4036
rect 4061 3904 4067 3916
rect 3981 3884 3987 3896
rect 4029 3864 4035 3876
rect 4093 3824 4099 3896
rect 4109 3884 4115 4136
rect 4157 4124 4163 4156
rect 4173 4144 4179 4276
rect 4269 4184 4275 4196
rect 4365 4143 4371 4256
rect 4381 4164 4387 4236
rect 4397 4204 4403 4316
rect 4413 4304 4419 4616
rect 4429 4324 4435 4576
rect 4525 4544 4531 4656
rect 4589 4604 4595 4636
rect 4637 4544 4643 4636
rect 4653 4584 4659 4656
rect 4717 4544 4723 4696
rect 4861 4664 4867 4716
rect 4909 4684 4915 4756
rect 4973 4664 4979 4736
rect 5005 4724 5011 4756
rect 4989 4704 4995 4716
rect 5021 4703 5027 4756
rect 5053 4724 5059 4756
rect 5165 4744 5171 4756
rect 5277 4724 5283 4736
rect 5037 4704 5043 4716
rect 5005 4697 5027 4703
rect 5005 4683 5011 4697
rect 4996 4677 5011 4683
rect 4749 4584 4755 4656
rect 4765 4564 4771 4616
rect 4621 4524 4627 4536
rect 4461 4384 4467 4436
rect 4413 4183 4419 4296
rect 4445 4184 4451 4316
rect 4413 4177 4435 4183
rect 4429 4164 4435 4177
rect 4324 4137 4355 4143
rect 4365 4137 4387 4143
rect 4349 4124 4355 4137
rect 4109 3744 4115 3876
rect 4173 3864 4179 3876
rect 4141 3844 4147 3856
rect 4205 3784 4211 3816
rect 4205 3764 4211 3776
rect 4077 3726 4083 3736
rect 3981 3644 3987 3716
rect 3933 3364 3939 3456
rect 3917 3344 3923 3356
rect 3860 3337 3884 3343
rect 3757 3324 3763 3336
rect 3965 3324 3971 3536
rect 3997 3484 4003 3496
rect 4109 3484 4115 3736
rect 3997 3384 4003 3396
rect 4013 3344 4019 3356
rect 4029 3344 4035 3456
rect 4060 3350 4068 3356
rect 4141 3344 4147 3496
rect 3725 3317 3740 3323
rect 3773 3303 3779 3316
rect 3661 3297 3779 3303
rect 3837 3284 3843 3316
rect 3981 3304 3987 3336
rect 4157 3324 4163 3376
rect 4173 3344 4179 3356
rect 4237 3344 4243 4096
rect 4269 3644 4275 3996
rect 4285 3764 4291 3796
rect 4301 3764 4307 4116
rect 4333 4104 4339 4116
rect 4317 4064 4323 4096
rect 4365 4084 4371 4116
rect 4317 4004 4323 4056
rect 4349 3984 4355 3996
rect 4381 3984 4387 4137
rect 4461 4084 4467 4336
rect 4477 4304 4483 4336
rect 4557 4304 4563 4476
rect 4637 4444 4643 4536
rect 4685 4504 4691 4516
rect 4717 4304 4723 4456
rect 4733 4444 4739 4556
rect 4781 4484 4787 4636
rect 4925 4524 4931 4656
rect 4973 4484 4979 4518
rect 4877 4464 4883 4476
rect 5005 4444 5011 4536
rect 5037 4524 5043 4656
rect 5069 4544 5075 4716
rect 5181 4704 5187 4716
rect 5101 4564 5107 4696
rect 5117 4684 5123 4696
rect 5133 4544 5139 4676
rect 5053 4504 5059 4536
rect 5133 4524 5139 4536
rect 5069 4484 5075 4516
rect 5165 4504 5171 4676
rect 5197 4644 5203 4716
rect 4509 4224 4515 4256
rect 4493 4164 4499 4196
rect 4509 4084 4515 4096
rect 4397 3963 4403 4036
rect 4477 4004 4483 4036
rect 4381 3957 4403 3963
rect 4365 3944 4371 3956
rect 4349 3923 4355 3936
rect 4349 3917 4371 3923
rect 4333 3844 4339 3896
rect 4365 3724 4371 3917
rect 4381 3904 4387 3957
rect 4397 3924 4403 3936
rect 4397 3764 4403 3796
rect 4429 3784 4435 3796
rect 4333 3644 4339 3696
rect 4253 3524 4259 3636
rect 4269 3563 4275 3636
rect 4269 3557 4291 3563
rect 4269 3524 4275 3536
rect 4205 3304 4211 3316
rect 4253 3304 4259 3516
rect 4285 3504 4291 3557
rect 4301 3364 4307 3596
rect 4317 3503 4323 3636
rect 4333 3604 4339 3636
rect 4381 3524 4387 3536
rect 4397 3504 4403 3716
rect 4445 3564 4451 3896
rect 4509 3584 4515 3894
rect 4525 3584 4531 4256
rect 4541 4144 4547 4156
rect 4557 4104 4563 4176
rect 4541 4024 4547 4076
rect 4573 3884 4579 4116
rect 4541 3784 4547 3836
rect 4621 3804 4627 4276
rect 4701 4244 4707 4296
rect 4781 4283 4787 4436
rect 4808 4406 4814 4414
rect 4822 4406 4828 4414
rect 4836 4406 4842 4414
rect 4850 4406 4856 4414
rect 4781 4277 4796 4283
rect 4701 4184 4707 4236
rect 4765 4184 4771 4216
rect 4781 4144 4787 4156
rect 4845 4144 4851 4196
rect 4861 4184 4867 4236
rect 4861 4164 4867 4176
rect 4877 4144 4883 4436
rect 4893 4304 4899 4316
rect 4925 4184 4931 4296
rect 4941 4224 4947 4336
rect 4957 4244 4963 4316
rect 4989 4304 4995 4416
rect 5133 4284 5139 4336
rect 5149 4284 5155 4316
rect 5181 4284 5187 4336
rect 4973 4264 4979 4276
rect 4940 4150 4948 4156
rect 4973 4144 4979 4176
rect 4685 4064 4691 4136
rect 4653 3924 4659 3936
rect 4669 3904 4675 3996
rect 4685 3844 4691 3936
rect 4557 3764 4563 3796
rect 4653 3744 4659 3756
rect 4669 3724 4675 3836
rect 4701 3784 4707 4136
rect 4717 3984 4723 4116
rect 4733 3944 4739 3956
rect 4733 3744 4739 3936
rect 4749 3904 4755 3996
rect 4781 3804 4787 4116
rect 4877 4024 4883 4056
rect 4808 4006 4814 4014
rect 4822 4006 4828 4014
rect 4836 4006 4842 4014
rect 4850 4006 4856 4014
rect 4893 3944 4899 4056
rect 4989 3944 4995 4276
rect 5021 4244 5027 4256
rect 5005 4144 5011 4196
rect 5021 4104 5027 4236
rect 5037 4124 5043 4156
rect 5053 4124 5059 4236
rect 5069 4204 5075 4236
rect 5085 4124 5091 4216
rect 5117 4164 5123 4196
rect 5149 4144 5155 4236
rect 5181 4184 5187 4276
rect 5213 4264 5219 4676
rect 5245 4564 5251 4596
rect 5261 4584 5267 4636
rect 5309 4564 5315 5056
rect 5501 5044 5507 5057
rect 5357 4904 5363 5036
rect 5517 4984 5523 4996
rect 5549 4984 5555 5016
rect 5533 4944 5539 4976
rect 5565 4944 5571 5076
rect 5597 5024 5603 5094
rect 5709 4984 5715 5236
rect 5837 5184 5843 5216
rect 5757 5064 5763 5076
rect 5741 4944 5747 5036
rect 5773 5004 5779 5076
rect 5789 5024 5795 5096
rect 5901 5064 5907 5356
rect 5997 5324 6003 5336
rect 6045 5324 6051 5376
rect 6221 5344 6227 5496
rect 6253 5484 6259 5496
rect 6253 5457 6268 5463
rect 6253 5344 6259 5457
rect 6285 5384 6291 5436
rect 6317 5383 6323 5496
rect 6381 5444 6387 5476
rect 6344 5406 6350 5414
rect 6358 5406 6364 5414
rect 6372 5406 6378 5414
rect 6386 5406 6392 5414
rect 6317 5377 6339 5383
rect 6317 5344 6323 5356
rect 5949 5124 5955 5176
rect 6029 5104 6035 5256
rect 6077 5104 6083 5316
rect 6141 5184 6147 5336
rect 6189 5243 6195 5276
rect 6173 5237 6195 5243
rect 6157 5163 6163 5236
rect 6173 5184 6179 5237
rect 6205 5204 6211 5316
rect 6141 5157 6163 5163
rect 6141 5124 6147 5157
rect 6205 5124 6211 5156
rect 5357 4724 5363 4896
rect 5373 4784 5379 4918
rect 5549 4884 5555 4896
rect 5453 4864 5459 4876
rect 5469 4864 5475 4876
rect 5341 4684 5347 4716
rect 5325 4664 5331 4676
rect 5389 4524 5395 4536
rect 5405 4504 5411 4836
rect 5437 4684 5443 4756
rect 5453 4684 5459 4716
rect 5453 4664 5459 4676
rect 5485 4664 5491 4716
rect 5501 4704 5507 4876
rect 5581 4864 5587 4916
rect 5549 4784 5555 4856
rect 5677 4784 5683 4916
rect 5693 4904 5699 4916
rect 5821 4784 5827 4856
rect 5517 4704 5523 4756
rect 5533 4684 5539 4716
rect 5597 4704 5603 4716
rect 5549 4664 5555 4696
rect 5661 4683 5667 4716
rect 5652 4677 5667 4683
rect 5501 4624 5507 4656
rect 5661 4584 5667 4677
rect 5693 4644 5699 4736
rect 5709 4584 5715 4656
rect 5757 4644 5763 4716
rect 5229 4304 5235 4396
rect 5293 4384 5299 4416
rect 5325 4384 5331 4476
rect 5421 4444 5427 4516
rect 5517 4484 5523 4536
rect 5629 4524 5635 4576
rect 5661 4544 5667 4576
rect 5693 4564 5699 4576
rect 5757 4564 5763 4636
rect 5773 4624 5779 4696
rect 5789 4664 5795 4676
rect 5677 4524 5683 4556
rect 5725 4544 5731 4556
rect 5757 4544 5763 4556
rect 5773 4544 5779 4596
rect 5789 4584 5795 4636
rect 5565 4484 5571 4496
rect 5613 4484 5619 4516
rect 5629 4504 5635 4516
rect 5725 4504 5731 4536
rect 5245 4264 5251 4276
rect 5309 4264 5315 4296
rect 5421 4284 5427 4436
rect 5805 4424 5811 4536
rect 5837 4524 5843 5036
rect 5869 4964 5875 5056
rect 5933 4926 5939 5076
rect 5997 4984 6003 5016
rect 6029 4944 6035 4956
rect 6061 4944 6067 5076
rect 6109 4924 6115 4936
rect 5965 4724 5971 4736
rect 5869 4604 5875 4636
rect 5885 4624 5891 4656
rect 5885 4544 5891 4556
rect 5837 4404 5843 4516
rect 5917 4504 5923 4636
rect 5933 4584 5939 4596
rect 5949 4584 5955 4656
rect 5997 4604 6003 4876
rect 6029 4704 6035 4776
rect 6045 4704 6051 4756
rect 6093 4564 6099 4716
rect 6141 4684 6147 5116
rect 6237 5104 6243 5136
rect 6269 5124 6275 5236
rect 6285 5104 6291 5336
rect 6333 5324 6339 5377
rect 6333 5284 6339 5296
rect 6333 5164 6339 5276
rect 6173 5084 6179 5096
rect 6157 5044 6163 5076
rect 6205 5063 6211 5096
rect 6221 5084 6227 5096
rect 6301 5084 6307 5156
rect 6349 5144 6355 5256
rect 6365 5184 6371 5376
rect 6381 5304 6387 5336
rect 6429 5304 6435 5436
rect 6349 5104 6355 5136
rect 6205 5057 6316 5063
rect 6381 5044 6387 5296
rect 6413 5124 6419 5136
rect 6429 5104 6435 5296
rect 6445 5264 6451 5316
rect 6461 5284 6467 5316
rect 6477 5304 6483 5476
rect 6557 5384 6563 5496
rect 6573 5484 6579 5496
rect 6589 5384 6595 5436
rect 6589 5344 6595 5356
rect 6573 5324 6579 5336
rect 6445 5204 6451 5236
rect 6461 5164 6467 5276
rect 6461 5124 6467 5156
rect 6525 5124 6531 5316
rect 6541 5264 6547 5296
rect 6541 5184 6547 5256
rect 6605 5164 6611 5496
rect 6621 5364 6627 5476
rect 6637 5384 6643 5476
rect 6653 5364 6659 5476
rect 6701 5464 6707 5536
rect 6781 5504 6787 5516
rect 6701 5384 6707 5436
rect 6717 5404 6723 5456
rect 6749 5444 6755 5496
rect 6797 5404 6803 5436
rect 6717 5344 6723 5396
rect 6733 5324 6739 5356
rect 6621 5304 6627 5316
rect 6701 5304 6707 5316
rect 6829 5224 6835 5496
rect 6909 5484 6915 5736
rect 6941 5684 6947 5696
rect 6957 5684 6963 5716
rect 7005 5704 7011 5716
rect 7021 5704 7027 5716
rect 6973 5664 6979 5696
rect 6989 5644 6995 5696
rect 6957 5504 6963 5636
rect 6909 5323 6915 5476
rect 7021 5324 7027 5336
rect 6909 5317 6924 5323
rect 6877 5304 6883 5316
rect 6493 5084 6499 5096
rect 6157 4864 6163 5036
rect 6344 5006 6350 5014
rect 6358 5006 6364 5014
rect 6372 5006 6378 5014
rect 6386 5006 6392 5014
rect 6285 4924 6291 4976
rect 6221 4884 6227 4916
rect 6205 4724 6211 4836
rect 6141 4644 6147 4656
rect 6157 4544 6163 4676
rect 6173 4644 6179 4696
rect 6205 4664 6211 4716
rect 6221 4684 6227 4856
rect 6317 4844 6323 4896
rect 6333 4784 6339 4936
rect 6413 4923 6419 5036
rect 6429 4924 6435 4936
rect 6404 4917 6419 4923
rect 6461 4744 6467 5076
rect 6525 5064 6531 5116
rect 6541 4924 6547 5076
rect 6237 4704 6243 4716
rect 6413 4684 6419 4716
rect 6461 4684 6467 4736
rect 6557 4724 6563 5056
rect 6573 5044 6579 5136
rect 6637 4964 6643 5036
rect 6701 5024 6707 5094
rect 6925 5084 6931 5316
rect 6989 5284 6995 5316
rect 7037 5084 7043 5436
rect 7053 5083 7059 5736
rect 7149 5724 7155 5736
rect 7197 5704 7203 5736
rect 7085 5544 7091 5696
rect 7101 5664 7107 5696
rect 7213 5684 7219 5716
rect 7133 5584 7139 5676
rect 7149 5544 7155 5676
rect 7117 5484 7123 5516
rect 7117 5464 7123 5476
rect 7085 5383 7091 5456
rect 7101 5404 7107 5436
rect 7069 5377 7091 5383
rect 7069 5344 7075 5377
rect 7133 5344 7139 5376
rect 7069 5084 7075 5116
rect 7053 5077 7068 5083
rect 7101 5083 7107 5296
rect 7117 5144 7123 5316
rect 7149 5284 7155 5536
rect 7165 5524 7171 5636
rect 7213 5584 7219 5656
rect 7229 5484 7235 5736
rect 7277 5584 7283 5636
rect 7325 5584 7331 5716
rect 7405 5584 7411 5636
rect 7325 5537 7340 5543
rect 7181 5343 7187 5456
rect 7245 5424 7251 5456
rect 7245 5344 7251 5396
rect 7261 5344 7267 5476
rect 7277 5384 7283 5496
rect 7325 5364 7331 5537
rect 7421 5504 7427 5536
rect 7341 5444 7347 5456
rect 7181 5337 7203 5343
rect 7165 5264 7171 5336
rect 7165 5164 7171 5236
rect 7133 5124 7139 5156
rect 7165 5104 7171 5136
rect 7101 5077 7116 5083
rect 6573 4784 6579 4836
rect 6589 4704 6595 4896
rect 6189 4543 6195 4636
rect 6269 4603 6275 4636
rect 6344 4606 6350 4614
rect 6358 4606 6364 4614
rect 6372 4606 6378 4614
rect 6386 4606 6392 4614
rect 6269 4597 6291 4603
rect 6285 4564 6291 4597
rect 6445 4584 6451 4676
rect 6477 4664 6483 4680
rect 6509 4644 6515 4656
rect 6525 4644 6531 4696
rect 6637 4684 6643 4956
rect 6653 4937 6668 4943
rect 6653 4904 6659 4937
rect 6733 4924 6739 5036
rect 6989 4984 6995 5016
rect 7005 4983 7011 5036
rect 7021 5024 7027 5056
rect 7005 4977 7027 4983
rect 6989 4957 7004 4963
rect 6733 4764 6739 4916
rect 6749 4884 6755 4936
rect 6685 4684 6691 4756
rect 6733 4724 6739 4736
rect 6797 4704 6803 4916
rect 6813 4724 6819 4956
rect 6813 4684 6819 4716
rect 6541 4664 6547 4676
rect 6573 4664 6579 4676
rect 6829 4664 6835 4756
rect 6845 4744 6851 4936
rect 6973 4924 6979 4936
rect 6957 4904 6963 4916
rect 6909 4884 6915 4896
rect 6925 4884 6931 4896
rect 6893 4764 6899 4876
rect 6925 4743 6931 4876
rect 6989 4784 6995 4957
rect 7021 4904 7027 4977
rect 7037 4964 7043 5076
rect 7197 5064 7203 5337
rect 7229 5284 7235 5316
rect 7325 5304 7331 5356
rect 7341 5324 7347 5436
rect 7389 5324 7395 5336
rect 7405 5324 7411 5376
rect 7421 5364 7427 5436
rect 7437 5303 7443 5736
rect 7453 5384 7459 5636
rect 7469 5504 7475 5516
rect 7437 5297 7459 5303
rect 7325 5243 7331 5296
rect 7325 5237 7347 5243
rect 7293 5104 7299 5156
rect 7341 5104 7347 5237
rect 7389 5144 7395 5236
rect 7213 5044 7219 5056
rect 7245 5044 7251 5096
rect 7293 5084 7299 5096
rect 7053 4984 7059 5036
rect 7133 4984 7139 5036
rect 7037 4924 7043 4936
rect 6916 4737 6931 4743
rect 6877 4664 6883 4736
rect 6909 4684 6915 4736
rect 7021 4724 7027 4896
rect 7085 4884 7091 4936
rect 6964 4717 6979 4723
rect 6973 4684 6979 4717
rect 7037 4704 7043 4716
rect 7053 4704 7059 4876
rect 7069 4704 7075 4756
rect 6989 4664 6995 4696
rect 7181 4684 7187 4936
rect 7277 4784 7283 5036
rect 7325 5024 7331 5096
rect 7373 4984 7379 5036
rect 7389 5004 7395 5056
rect 7405 5024 7411 5056
rect 7421 5024 7427 5056
rect 7405 4983 7411 5016
rect 7380 4977 7395 4983
rect 7405 4977 7420 4983
rect 7389 4964 7395 4977
rect 7405 4763 7411 4836
rect 7405 4757 7427 4763
rect 7293 4704 7299 4716
rect 7405 4704 7411 4736
rect 7421 4684 7427 4757
rect 6621 4564 6627 4576
rect 6781 4564 6787 4636
rect 6493 4544 6499 4556
rect 6525 4544 6531 4556
rect 6180 4537 6195 4543
rect 5757 4344 5763 4356
rect 5869 4344 5875 4436
rect 5469 4304 5475 4336
rect 5245 4184 5251 4216
rect 5325 4184 5331 4196
rect 5229 4164 5235 4176
rect 5341 4164 5347 4276
rect 4557 3704 4563 3718
rect 4605 3644 4611 3676
rect 4621 3584 4627 3716
rect 4781 3704 4787 3716
rect 4637 3584 4643 3696
rect 4813 3644 4819 3736
rect 4829 3724 4835 3756
rect 4861 3664 4867 3876
rect 4941 3844 4947 3896
rect 4685 3564 4691 3636
rect 4808 3606 4814 3614
rect 4822 3606 4828 3614
rect 4836 3606 4842 3614
rect 4850 3606 4856 3614
rect 4509 3523 4515 3536
rect 4749 3524 4755 3596
rect 4509 3517 4547 3523
rect 4445 3504 4451 3516
rect 4317 3497 4332 3503
rect 4301 3344 4307 3356
rect 4333 3344 4339 3456
rect 4365 3424 4371 3456
rect 4397 3384 4403 3496
rect 4493 3484 4499 3516
rect 4541 3503 4547 3517
rect 4621 3504 4627 3516
rect 4541 3497 4556 3503
rect 4429 3444 4435 3476
rect 4477 3364 4483 3476
rect 3645 3124 3651 3136
rect 3565 3104 3571 3116
rect 3421 3097 3443 3103
rect 3421 3084 3427 3097
rect 3652 3097 3676 3103
rect 3453 3084 3459 3096
rect 3245 3037 3267 3043
rect 2493 2644 2499 2676
rect 2637 2644 2643 2656
rect 2525 2584 2531 2616
rect 2557 2584 2563 2636
rect 2669 2624 2675 2696
rect 2733 2664 2739 2694
rect 2797 2684 2803 2696
rect 2653 2564 2659 2596
rect 2797 2564 2803 2676
rect 2573 2544 2579 2556
rect 2861 2544 2867 2596
rect 2877 2564 2883 2636
rect 2909 2584 2915 2696
rect 3021 2684 3027 2936
rect 3197 2844 3203 2956
rect 3245 2784 3251 3037
rect 3272 3006 3278 3014
rect 3286 3006 3292 3014
rect 3300 3006 3306 3014
rect 3314 3006 3320 3014
rect 3341 2944 3347 3056
rect 3437 2984 3443 3076
rect 3373 2944 3379 2976
rect 3453 2924 3459 2956
rect 3325 2884 3331 2916
rect 3469 2904 3475 2996
rect 3517 2984 3523 3056
rect 3533 3004 3539 3096
rect 3693 3084 3699 3136
rect 3789 3104 3795 3156
rect 3917 3144 3923 3296
rect 4205 3204 4211 3256
rect 3789 3084 3795 3096
rect 3597 3077 3612 3083
rect 3549 3064 3555 3076
rect 3501 2944 3507 2976
rect 3517 2944 3523 2976
rect 3533 2964 3539 2976
rect 3549 2964 3555 3016
rect 3565 2984 3571 3076
rect 3597 2984 3603 3077
rect 3677 2984 3683 3076
rect 3725 2984 3731 3056
rect 3773 3024 3779 3076
rect 3805 3064 3811 3076
rect 3885 3064 3891 3136
rect 3981 3104 3987 3116
rect 4205 3084 4211 3196
rect 4253 3184 4259 3236
rect 3485 2883 3491 2936
rect 3549 2884 3555 2956
rect 3645 2944 3651 2976
rect 3661 2944 3667 2956
rect 3757 2944 3763 2976
rect 3773 2944 3779 2956
rect 3837 2944 3843 3056
rect 3565 2937 3603 2943
rect 3485 2877 3523 2883
rect 3517 2863 3523 2877
rect 3565 2863 3571 2937
rect 3581 2864 3587 2916
rect 3597 2904 3603 2937
rect 3805 2904 3811 2936
rect 3869 2924 3875 3036
rect 3885 2964 3891 3016
rect 3901 2984 3907 2996
rect 3517 2857 3571 2863
rect 3117 2664 3123 2776
rect 3245 2744 3251 2776
rect 3165 2664 3171 2696
rect 3485 2684 3491 2696
rect 2957 2584 2963 2636
rect 2973 2544 2979 2596
rect 3085 2544 3091 2576
rect 3101 2564 3107 2596
rect 3197 2584 3203 2656
rect 3245 2584 3251 2656
rect 3272 2606 3278 2614
rect 3286 2606 3292 2614
rect 3300 2606 3306 2614
rect 3314 2606 3320 2614
rect 2429 2504 2435 2516
rect 2461 2304 2467 2376
rect 2477 2284 2483 2536
rect 2909 2524 2915 2536
rect 2637 2364 2643 2436
rect 2621 2304 2627 2316
rect 2669 2304 2675 2436
rect 2685 2384 2691 2496
rect 2797 2464 2803 2518
rect 2989 2504 2995 2516
rect 2957 2484 2963 2496
rect 2925 2324 2931 2356
rect 3021 2344 3027 2536
rect 3149 2523 3155 2556
rect 3149 2517 3164 2523
rect 3037 2504 3043 2516
rect 3181 2504 3187 2536
rect 3229 2524 3235 2556
rect 3245 2504 3251 2576
rect 3261 2524 3267 2556
rect 3357 2504 3363 2536
rect 3357 2484 3363 2496
rect 3053 2384 3059 2456
rect 2724 2297 2739 2303
rect 2573 2244 2579 2256
rect 2589 2244 2595 2276
rect 2637 2264 2643 2296
rect 2573 2184 2579 2216
rect 2317 1884 2323 1936
rect 2381 1903 2387 2136
rect 2429 2124 2435 2176
rect 2541 2143 2547 2176
rect 2541 2137 2556 2143
rect 2557 2124 2563 2136
rect 2573 2084 2579 2136
rect 2589 2124 2595 2236
rect 2621 2204 2627 2236
rect 2637 2163 2643 2236
rect 2653 2224 2659 2276
rect 2685 2204 2691 2276
rect 2708 2257 2716 2263
rect 2621 2157 2643 2163
rect 2605 2103 2611 2136
rect 2621 2124 2627 2157
rect 2605 2097 2627 2103
rect 2621 1984 2627 2097
rect 2637 1984 2643 2136
rect 2653 2124 2659 2196
rect 2701 2164 2707 2256
rect 2733 2164 2739 2297
rect 2916 2297 2931 2303
rect 2765 2164 2771 2296
rect 2797 2224 2803 2296
rect 2701 2004 2707 2156
rect 2733 2124 2739 2156
rect 2765 2144 2771 2156
rect 2797 2144 2803 2216
rect 2813 2184 2819 2236
rect 2861 2184 2867 2196
rect 2925 2184 2931 2297
rect 2989 2284 2995 2316
rect 3005 2304 3011 2316
rect 3149 2304 3155 2316
rect 2957 2264 2963 2276
rect 3005 2184 3011 2296
rect 3101 2284 3107 2296
rect 2845 2144 2851 2176
rect 3037 2164 3043 2276
rect 3085 2184 3091 2276
rect 3117 2183 3123 2236
rect 3149 2184 3155 2276
rect 3181 2184 3187 2396
rect 3197 2384 3203 2476
rect 3229 2317 3244 2323
rect 3229 2304 3235 2317
rect 3261 2304 3267 2436
rect 3373 2284 3379 2676
rect 3389 2544 3395 2656
rect 3421 2564 3427 2656
rect 3453 2644 3459 2656
rect 3453 2584 3459 2616
rect 3437 2524 3443 2556
rect 3469 2524 3475 2556
rect 3501 2544 3507 2676
rect 3469 2484 3475 2516
rect 3485 2504 3491 2536
rect 3501 2524 3507 2536
rect 3272 2206 3278 2214
rect 3286 2206 3292 2214
rect 3300 2206 3306 2214
rect 3314 2206 3320 2214
rect 3117 2177 3139 2183
rect 3021 2144 3027 2156
rect 3068 2150 3076 2156
rect 3133 2144 3139 2177
rect 3165 2164 3171 2176
rect 3341 2144 3347 2276
rect 3501 2184 3507 2236
rect 3517 2144 3523 2836
rect 3885 2744 3891 2956
rect 3981 2944 3987 2956
rect 3997 2924 4003 2936
rect 3933 2844 3939 2916
rect 4045 2904 4051 2996
rect 4205 2943 4211 3076
rect 4189 2937 4211 2943
rect 3949 2884 3955 2896
rect 4077 2864 4083 2916
rect 3549 2724 3555 2736
rect 3533 2717 3548 2723
rect 3533 2664 3539 2717
rect 3597 2664 3603 2676
rect 3533 2504 3539 2576
rect 3565 2523 3571 2636
rect 3565 2517 3580 2523
rect 3661 2484 3667 2518
rect 3533 2384 3539 2476
rect 3693 2384 3699 2656
rect 3709 2584 3715 2696
rect 3789 2684 3795 2736
rect 3837 2684 3843 2716
rect 3965 2704 3971 2836
rect 4093 2784 4099 2936
rect 3853 2677 3868 2683
rect 3725 2624 3731 2676
rect 3757 2664 3763 2676
rect 3837 2584 3843 2656
rect 3821 2544 3827 2556
rect 3709 2304 3715 2516
rect 3725 2284 3731 2296
rect 3757 2284 3763 2296
rect 3533 2224 3539 2236
rect 3677 2144 3683 2276
rect 2749 2104 2755 2136
rect 2893 2124 2899 2136
rect 2925 2124 2931 2136
rect 3021 2124 3027 2136
rect 2765 2104 2771 2116
rect 2781 2084 2787 2116
rect 2893 2104 2899 2116
rect 2861 2084 2867 2096
rect 2445 1924 2451 1936
rect 2365 1897 2387 1903
rect 2365 1744 2371 1897
rect 2493 1884 2499 1956
rect 2525 1864 2531 1876
rect 2557 1864 2563 1956
rect 2669 1884 2675 1916
rect 2749 1884 2755 1916
rect 2589 1864 2595 1880
rect 2509 1784 2515 1836
rect 2541 1804 2547 1836
rect 2429 1744 2435 1776
rect 2557 1744 2563 1856
rect 2605 1784 2611 1816
rect 2333 1704 2339 1718
rect 2349 1584 2355 1636
rect 2365 1543 2371 1736
rect 2365 1537 2387 1543
rect 2173 1404 2179 1476
rect 2189 1363 2195 1436
rect 2221 1364 2227 1476
rect 2253 1424 2259 1516
rect 2301 1484 2307 1496
rect 2381 1484 2387 1537
rect 2413 1502 2419 1716
rect 2445 1684 2451 1716
rect 2461 1644 2467 1736
rect 2557 1703 2563 1736
rect 2589 1724 2595 1776
rect 2685 1764 2691 1876
rect 2701 1864 2707 1876
rect 2637 1744 2643 1756
rect 2557 1697 2572 1703
rect 2685 1664 2691 1756
rect 2717 1724 2723 1756
rect 2733 1704 2739 1836
rect 2765 1744 2771 1996
rect 2797 1884 2803 1956
rect 2813 1884 2819 2056
rect 2829 1904 2835 1976
rect 2877 1864 2883 1976
rect 2973 1904 2979 1936
rect 3165 1924 3171 2096
rect 3005 1864 3011 1876
rect 2781 1784 2787 1816
rect 2541 1584 2547 1656
rect 2589 1484 2595 1576
rect 2669 1504 2675 1516
rect 2269 1444 2275 1456
rect 2301 1364 2307 1416
rect 2621 1364 2627 1476
rect 2109 1357 2131 1363
rect 2029 1164 2035 1336
rect 2061 1304 2067 1356
rect 2125 1344 2131 1357
rect 2173 1357 2195 1363
rect 2045 1204 2051 1236
rect 2013 984 2019 1036
rect 1933 924 1939 936
rect 1981 904 1987 936
rect 1981 704 1987 896
rect 2045 784 2051 1056
rect 2061 1044 2067 1296
rect 2109 1084 2115 1336
rect 2157 1304 2163 1336
rect 2173 1324 2179 1357
rect 2237 1284 2243 1316
rect 2125 1144 2131 1276
rect 2221 1224 2227 1236
rect 2141 1104 2147 1196
rect 2157 1084 2163 1096
rect 2301 1084 2307 1356
rect 2317 1124 2323 1156
rect 2333 1084 2339 1136
rect 2349 1084 2355 1236
rect 2365 1144 2371 1336
rect 2397 1204 2403 1296
rect 2397 1164 2403 1196
rect 2413 1124 2419 1176
rect 2429 1124 2435 1236
rect 2461 1184 2467 1336
rect 2685 1324 2691 1636
rect 2749 1624 2755 1696
rect 2765 1584 2771 1736
rect 2813 1724 2819 1856
rect 2829 1744 2835 1796
rect 2781 1584 2787 1636
rect 2797 1584 2803 1696
rect 2861 1604 2867 1836
rect 2893 1824 2899 1836
rect 2877 1724 2883 1776
rect 2893 1684 2899 1696
rect 2909 1504 2915 1836
rect 2941 1744 2947 1796
rect 2957 1684 2963 1716
rect 2989 1644 2995 1676
rect 3005 1524 3011 1736
rect 3021 1684 3027 1896
rect 3037 1884 3043 1896
rect 3069 1864 3075 1916
rect 3181 1904 3187 2036
rect 3229 1924 3235 1936
rect 3085 1864 3091 1896
rect 3133 1884 3139 1896
rect 3181 1864 3187 1876
rect 3213 1844 3219 1916
rect 3261 1884 3267 1896
rect 3277 1884 3283 2016
rect 3357 1964 3363 2076
rect 3373 1984 3379 2076
rect 3437 1984 3443 2116
rect 3245 1784 3251 1816
rect 3272 1806 3278 1814
rect 3286 1806 3292 1814
rect 3300 1806 3306 1814
rect 3314 1806 3320 1814
rect 3037 1724 3043 1756
rect 3053 1744 3059 1756
rect 3069 1724 3075 1776
rect 3101 1724 3107 1756
rect 3213 1744 3219 1756
rect 3277 1744 3283 1756
rect 3325 1744 3331 1776
rect 3357 1764 3363 1956
rect 3373 1844 3379 1896
rect 3389 1864 3395 1876
rect 3373 1764 3379 1836
rect 3421 1744 3427 1936
rect 3453 1924 3459 2016
rect 3437 1884 3443 1896
rect 3437 1784 3443 1876
rect 3453 1804 3459 1916
rect 3469 1864 3475 1956
rect 3453 1743 3459 1796
rect 3444 1737 3459 1743
rect 3021 1584 3027 1656
rect 3117 1644 3123 1716
rect 3149 1704 3155 1736
rect 3165 1704 3171 1736
rect 3181 1724 3187 1736
rect 3261 1724 3267 1736
rect 3357 1724 3363 1736
rect 3412 1717 3436 1723
rect 3261 1704 3267 1716
rect 3405 1664 3411 1696
rect 3453 1644 3459 1676
rect 3133 1624 3139 1636
rect 3213 1584 3219 1636
rect 3261 1504 3267 1536
rect 3357 1504 3363 1636
rect 3469 1504 3475 1856
rect 2717 1484 2723 1496
rect 3421 1484 3427 1494
rect 2477 1144 2483 1156
rect 2397 1084 2403 1116
rect 2493 1104 2499 1316
rect 2621 1284 2627 1318
rect 2509 1124 2515 1136
rect 2573 1124 2579 1236
rect 2077 1024 2083 1056
rect 2301 1044 2307 1076
rect 2333 1064 2339 1076
rect 2381 1064 2387 1076
rect 2445 1044 2451 1076
rect 2125 904 2131 936
rect 2173 924 2179 1036
rect 2205 944 2211 976
rect 2221 924 2227 996
rect 2253 984 2259 1036
rect 2461 964 2467 996
rect 2525 964 2531 1016
rect 2061 684 2067 816
rect 2173 784 2179 896
rect 2269 744 2275 836
rect 2397 784 2403 918
rect 1677 584 1683 616
rect 1885 603 1891 676
rect 2061 604 2067 676
rect 2205 664 2211 736
rect 1869 597 1891 603
rect 1524 577 1539 583
rect 1229 477 1251 483
rect 1229 384 1235 456
rect 1245 304 1251 477
rect 1389 443 1395 536
rect 1405 524 1411 576
rect 1869 564 1875 597
rect 2253 584 2259 696
rect 2333 684 2339 696
rect 2349 684 2355 756
rect 2381 724 2387 736
rect 2477 724 2483 836
rect 2381 697 2396 703
rect 1645 544 1651 556
rect 1869 526 1875 536
rect 1645 504 1651 516
rect 1373 437 1395 443
rect 1309 324 1315 436
rect 1373 284 1379 437
rect 1736 406 1742 414
rect 1750 406 1756 414
rect 1764 406 1770 414
rect 1778 406 1784 414
rect 1837 384 1843 516
rect 1565 344 1571 356
rect 1421 304 1427 336
rect 1037 124 1043 276
rect 1165 184 1171 256
rect 1373 243 1379 276
rect 1357 237 1379 243
rect 1309 224 1315 236
rect 1181 177 1196 183
rect 1181 144 1187 177
rect 1197 164 1203 176
rect 1357 144 1363 237
rect 1389 144 1395 216
rect 1053 124 1059 136
rect 1149 124 1155 136
rect 356 97 371 103
rect 205 84 211 96
rect 941 84 947 96
rect 957 84 963 116
rect 1389 84 1395 116
rect 1453 104 1459 316
rect 1501 144 1507 256
rect 1565 184 1571 296
rect 1613 244 1619 256
rect 1677 243 1683 296
rect 1693 264 1699 276
rect 1677 237 1699 243
rect 1629 184 1635 216
rect 1693 184 1699 237
rect 1533 143 1539 156
rect 1613 144 1619 156
rect 1677 144 1683 156
rect 1517 137 1539 143
rect 1517 124 1523 137
rect 1613 104 1619 136
rect 1693 124 1699 176
rect 1725 144 1731 256
rect 1741 224 1747 296
rect 1757 284 1763 316
rect 1901 304 1907 536
rect 1933 484 1939 556
rect 2125 544 2131 556
rect 2253 524 2259 576
rect 2269 544 2275 676
rect 2285 624 2291 636
rect 2285 540 2291 616
rect 2317 584 2323 656
rect 2349 564 2355 676
rect 2381 584 2387 697
rect 2429 684 2435 696
rect 2493 684 2499 756
rect 2541 744 2547 936
rect 2589 903 2595 1216
rect 2605 1103 2611 1176
rect 2605 1097 2620 1103
rect 2637 1084 2643 1236
rect 2669 1184 2675 1276
rect 2653 1104 2659 1116
rect 2637 1044 2643 1076
rect 2669 1064 2675 1096
rect 2717 1084 2723 1236
rect 2797 1224 2803 1436
rect 2861 1344 2867 1476
rect 3357 1444 3363 1456
rect 3272 1406 3278 1414
rect 3286 1406 3292 1414
rect 3300 1406 3306 1414
rect 3314 1406 3320 1414
rect 3389 1384 3395 1476
rect 2909 1364 2915 1376
rect 3069 1304 3075 1336
rect 3117 1284 3123 1316
rect 3213 1304 3219 1336
rect 3389 1304 3395 1376
rect 3485 1303 3491 2076
rect 3501 1984 3507 2096
rect 3533 2084 3539 2136
rect 3629 2104 3635 2136
rect 3661 2124 3667 2136
rect 3645 2004 3651 2116
rect 3661 1904 3667 2016
rect 3693 1904 3699 2036
rect 3709 1964 3715 2156
rect 3757 2024 3763 2276
rect 3821 2264 3827 2536
rect 3853 2224 3859 2677
rect 3901 2524 3907 2676
rect 3901 2343 3907 2436
rect 3933 2384 3939 2536
rect 4013 2524 4019 2616
rect 4077 2584 4083 2676
rect 4109 2604 4115 2896
rect 4125 2864 4131 2916
rect 4141 2884 4147 2916
rect 4189 2683 4195 2937
rect 4285 2924 4291 2956
rect 4205 2784 4211 2916
rect 4301 2824 4307 3096
rect 4317 2944 4323 3236
rect 4333 3064 4339 3336
rect 4365 2884 4371 3316
rect 4365 2864 4371 2876
rect 4237 2704 4243 2756
rect 4189 2677 4204 2683
rect 4029 2564 4035 2576
rect 4093 2544 4099 2596
rect 4173 2584 4179 2676
rect 4189 2564 4195 2677
rect 4269 2624 4275 2636
rect 4317 2624 4323 2716
rect 4365 2684 4371 2796
rect 4381 2684 4387 3236
rect 4493 3184 4499 3476
rect 4509 3184 4515 3496
rect 4525 3244 4531 3318
rect 4557 3184 4563 3476
rect 4589 3364 4595 3496
rect 4605 3384 4611 3496
rect 4701 3484 4707 3496
rect 4621 3384 4627 3476
rect 4669 3424 4675 3476
rect 4749 3464 4755 3516
rect 4829 3504 4835 3516
rect 4797 3484 4803 3496
rect 4797 3464 4803 3476
rect 4685 3384 4691 3396
rect 4605 3324 4611 3376
rect 4717 3344 4723 3356
rect 4749 3344 4755 3396
rect 4797 3384 4803 3436
rect 4829 3384 4835 3416
rect 4781 3324 4787 3356
rect 4813 3344 4819 3356
rect 4733 3284 4739 3316
rect 4808 3206 4814 3214
rect 4822 3206 4828 3214
rect 4836 3206 4842 3214
rect 4850 3206 4856 3214
rect 4877 3184 4883 3816
rect 4957 3764 4963 3836
rect 4973 3824 4979 3856
rect 4989 3744 4995 3876
rect 5053 3764 5059 3816
rect 4909 3664 4915 3716
rect 4957 3504 4963 3516
rect 4909 3444 4915 3476
rect 4973 3444 4979 3516
rect 4957 3384 4963 3436
rect 4900 3340 4915 3343
rect 4900 3337 4908 3340
rect 4893 3184 4899 3336
rect 4973 3304 4979 3316
rect 4989 3264 4995 3736
rect 5021 3664 5027 3716
rect 5085 3544 5091 4076
rect 5165 3883 5171 3936
rect 5197 3924 5203 4096
rect 5213 4024 5219 4136
rect 5229 4024 5235 4156
rect 5293 4124 5299 4136
rect 5277 4004 5283 4116
rect 5309 4104 5315 4156
rect 5357 4144 5363 4280
rect 5373 4124 5379 4136
rect 5389 4124 5395 4236
rect 5453 4144 5459 4196
rect 5229 3984 5235 3996
rect 5181 3917 5196 3923
rect 5181 3904 5187 3917
rect 5261 3904 5267 3936
rect 5325 3924 5331 4036
rect 5357 3984 5363 4116
rect 5373 4064 5379 4116
rect 5453 3924 5459 3956
rect 5485 3944 5491 4136
rect 5156 3880 5171 3883
rect 5149 3877 5171 3880
rect 5101 3764 5107 3836
rect 5181 3584 5187 3896
rect 5293 3864 5299 3876
rect 5309 3764 5315 3876
rect 5325 3764 5331 3896
rect 5405 3884 5411 3896
rect 5501 3884 5507 4296
rect 5549 4184 5555 4276
rect 5597 4244 5603 4276
rect 5661 4264 5667 4296
rect 5709 4284 5715 4296
rect 5597 4184 5603 4216
rect 5517 4144 5523 4156
rect 5517 3924 5523 4116
rect 5565 4104 5571 4136
rect 5613 4104 5619 4116
rect 5661 4104 5667 4156
rect 5693 4144 5699 4156
rect 5725 4104 5731 4296
rect 5741 4164 5747 4336
rect 5757 4184 5763 4276
rect 5789 4184 5795 4256
rect 5821 4224 5827 4296
rect 5869 4284 5875 4336
rect 5885 4304 5891 4356
rect 5837 4244 5843 4276
rect 5901 4264 5907 4296
rect 5933 4264 5939 4436
rect 6029 4324 6035 4336
rect 5997 4264 6003 4296
rect 5853 4204 5859 4236
rect 5933 4224 5939 4256
rect 5757 4143 5763 4156
rect 5748 4137 5763 4143
rect 5773 4124 5779 4156
rect 5821 4144 5827 4156
rect 5853 4144 5859 4176
rect 5869 4144 5875 4216
rect 5869 4124 5875 4136
rect 6013 4126 6019 4156
rect 6045 4144 6051 4536
rect 6061 4484 6067 4518
rect 6541 4524 6547 4536
rect 6701 4524 6707 4556
rect 6205 4504 6211 4516
rect 6221 4504 6227 4516
rect 6285 4504 6291 4518
rect 6637 4517 6652 4523
rect 6109 4384 6115 4476
rect 6125 4464 6131 4496
rect 6413 4484 6419 4496
rect 6477 4384 6483 4516
rect 6605 4384 6611 4516
rect 6637 4384 6643 4517
rect 6653 4504 6659 4516
rect 6669 4484 6675 4496
rect 6749 4484 6755 4556
rect 6781 4544 6787 4556
rect 6797 4524 6803 4576
rect 6749 4444 6755 4476
rect 6157 4324 6163 4336
rect 6205 4324 6211 4336
rect 6077 4184 6083 4296
rect 6100 4277 6115 4283
rect 6109 4156 6115 4277
rect 6141 4264 6147 4296
rect 6173 4284 6179 4316
rect 6237 4304 6243 4316
rect 6141 4184 6147 4216
rect 6173 4144 6179 4276
rect 6189 4244 6195 4296
rect 6253 4224 6259 4276
rect 6285 4264 6291 4316
rect 6301 4284 6307 4356
rect 6381 4304 6387 4316
rect 6317 4264 6323 4296
rect 6461 4263 6467 4316
rect 6605 4304 6611 4376
rect 6797 4344 6803 4516
rect 6685 4284 6691 4336
rect 6493 4264 6499 4276
rect 6445 4257 6467 4263
rect 6077 4124 6083 4136
rect 5613 3984 5619 3996
rect 5261 3584 5267 3718
rect 5405 3704 5411 3876
rect 5421 3783 5427 3856
rect 5533 3784 5539 3896
rect 5629 3884 5635 4016
rect 5661 4004 5667 4096
rect 5821 4024 5827 4056
rect 5821 3924 5827 4016
rect 5837 3924 5843 4116
rect 5885 4004 5891 4036
rect 5853 3944 5859 3956
rect 5693 3884 5699 3896
rect 5629 3864 5635 3876
rect 5757 3864 5763 3896
rect 5789 3884 5795 3896
rect 5821 3864 5827 3916
rect 5853 3864 5859 3896
rect 5901 3884 5907 3916
rect 5933 3884 5939 3896
rect 5997 3864 6003 3896
rect 5789 3784 5795 3816
rect 5869 3784 5875 3796
rect 5421 3777 5443 3783
rect 5437 3744 5443 3777
rect 5821 3757 5836 3763
rect 5293 3564 5299 3656
rect 5437 3624 5443 3736
rect 5501 3604 5507 3716
rect 5437 3584 5443 3596
rect 5405 3537 5523 3543
rect 5037 3484 5043 3496
rect 5005 3384 5011 3476
rect 5005 3364 5011 3376
rect 5021 3364 5027 3436
rect 5021 3323 5027 3356
rect 5021 3317 5036 3323
rect 5053 3284 5059 3436
rect 5069 3263 5075 3436
rect 5085 3344 5091 3456
rect 5197 3424 5203 3476
rect 5213 3464 5219 3496
rect 5229 3484 5235 3496
rect 5261 3464 5267 3516
rect 5277 3464 5283 3476
rect 5325 3464 5331 3536
rect 5373 3524 5379 3536
rect 5405 3524 5411 3537
rect 5517 3524 5523 3537
rect 5341 3464 5347 3496
rect 5325 3404 5331 3456
rect 5357 3424 5363 3516
rect 5373 3484 5379 3516
rect 5421 3504 5427 3516
rect 5501 3504 5507 3516
rect 5405 3484 5411 3496
rect 5421 3464 5427 3496
rect 5437 3443 5443 3476
rect 5421 3437 5443 3443
rect 5101 3324 5107 3376
rect 5133 3304 5139 3316
rect 5181 3304 5187 3376
rect 5261 3364 5267 3396
rect 5229 3324 5235 3336
rect 5069 3257 5091 3263
rect 5053 3184 5059 3236
rect 4413 3064 4419 3116
rect 4445 3064 4451 3076
rect 4397 3024 4403 3036
rect 4429 2924 4435 2936
rect 4445 2924 4451 3056
rect 4397 2884 4403 2896
rect 4413 2704 4419 2716
rect 4445 2704 4451 2896
rect 4461 2684 4467 2916
rect 4493 2903 4499 3136
rect 4509 3104 4515 3136
rect 4605 3124 4611 3156
rect 4525 2944 4531 3056
rect 4541 3044 4547 3076
rect 4557 3064 4563 3096
rect 4541 2964 4547 3016
rect 4509 2904 4515 2916
rect 4541 2904 4547 2956
rect 4573 2944 4579 3116
rect 4637 3104 4643 3136
rect 4653 3084 4659 3116
rect 4637 3044 4643 3056
rect 4669 3044 4675 3116
rect 4637 2944 4643 3036
rect 4685 2924 4691 3136
rect 4717 3084 4723 3156
rect 4765 3124 4771 3176
rect 4733 2944 4739 3116
rect 5069 3104 5075 3236
rect 4996 3097 5011 3103
rect 4749 2964 4755 3076
rect 4493 2897 4508 2903
rect 4541 2804 4547 2896
rect 4685 2844 4691 2916
rect 4573 2784 4579 2836
rect 4669 2764 4675 2836
rect 4749 2824 4755 2836
rect 4509 2684 4515 2736
rect 4205 2544 4211 2576
rect 4301 2564 4307 2576
rect 4109 2504 4115 2516
rect 3901 2337 3923 2343
rect 3773 2164 3779 2196
rect 3837 2144 3843 2156
rect 3757 1964 3763 1996
rect 3789 1924 3795 2076
rect 3821 1964 3827 2116
rect 3821 1944 3827 1956
rect 3837 1924 3843 2096
rect 3853 2084 3859 2136
rect 3901 2104 3907 2156
rect 3533 1824 3539 1856
rect 3597 1764 3603 1896
rect 3773 1804 3779 1856
rect 3501 1744 3507 1756
rect 3597 1744 3603 1756
rect 3501 1684 3507 1716
rect 3517 1644 3523 1716
rect 3533 1524 3539 1636
rect 3565 1604 3571 1736
rect 3629 1724 3635 1776
rect 3645 1764 3651 1796
rect 3741 1744 3747 1796
rect 3821 1764 3827 1856
rect 3853 1804 3859 2076
rect 3901 1944 3907 1956
rect 3885 1884 3891 1896
rect 3917 1884 3923 2337
rect 3965 2284 3971 2296
rect 3933 2004 3939 2116
rect 3965 2024 3971 2276
rect 3981 2184 3987 2316
rect 4013 2184 4019 2296
rect 4061 2264 4067 2296
rect 4077 2284 4083 2376
rect 4029 2104 4035 2136
rect 4109 2124 4115 2456
rect 4237 2344 4243 2436
rect 4253 2364 4259 2516
rect 4269 2484 4275 2516
rect 4301 2384 4307 2556
rect 4317 2424 4323 2616
rect 4349 2464 4355 2496
rect 4365 2444 4371 2676
rect 4461 2664 4467 2676
rect 4477 2584 4483 2616
rect 4541 2584 4547 2716
rect 4621 2704 4627 2736
rect 4781 2724 4787 3056
rect 4909 3024 4915 3096
rect 4957 2944 4963 3076
rect 4973 3064 4979 3076
rect 4973 2984 4979 3016
rect 5005 2924 5011 3097
rect 5069 3044 5075 3056
rect 5085 2944 5091 3257
rect 5101 3144 5107 3236
rect 5165 3144 5171 3296
rect 5165 2984 5171 3136
rect 5197 3124 5203 3296
rect 5261 3184 5267 3356
rect 5325 3324 5331 3356
rect 5357 3344 5363 3376
rect 5197 3084 5203 3094
rect 5341 3084 5347 3336
rect 5389 3304 5395 3436
rect 5405 3344 5411 3416
rect 5421 3384 5427 3437
rect 5437 3364 5443 3396
rect 5453 3364 5459 3496
rect 5469 3444 5475 3476
rect 5437 3304 5443 3356
rect 5485 3324 5491 3456
rect 5501 3424 5507 3476
rect 5517 3464 5523 3496
rect 5533 3384 5539 3696
rect 5677 3664 5683 3718
rect 5581 3464 5587 3636
rect 5668 3517 5683 3523
rect 5620 3497 5644 3503
rect 5677 3503 5683 3517
rect 5677 3497 5692 3503
rect 5677 3444 5683 3497
rect 5581 3364 5587 3376
rect 5517 3303 5523 3336
rect 5501 3297 5523 3303
rect 5501 3184 5507 3297
rect 5565 3284 5571 3316
rect 5613 3304 5619 3376
rect 5661 3364 5667 3416
rect 5677 3384 5683 3436
rect 5709 3384 5715 3736
rect 5789 3724 5795 3736
rect 5741 3684 5747 3716
rect 5821 3704 5827 3757
rect 5837 3704 5843 3736
rect 5789 3584 5795 3656
rect 5757 3504 5763 3516
rect 5789 3504 5795 3556
rect 5821 3464 5827 3696
rect 5668 3357 5683 3363
rect 5677 3184 5683 3357
rect 5709 3324 5715 3356
rect 5773 3144 5779 3456
rect 5837 3424 5843 3456
rect 5805 3263 5811 3336
rect 5805 3257 5827 3263
rect 5821 3184 5827 3257
rect 5853 3184 5859 3416
rect 5885 3384 5891 3836
rect 5917 3724 5923 3736
rect 5901 3544 5907 3716
rect 5917 3664 5923 3716
rect 5933 3704 5939 3796
rect 6029 3784 6035 3896
rect 6061 3844 6067 3856
rect 6077 3804 6083 4116
rect 6205 3924 6211 4196
rect 6269 4164 6275 4236
rect 6344 4206 6350 4214
rect 6358 4206 6364 4214
rect 6372 4206 6378 4214
rect 6386 4206 6392 4214
rect 6317 4126 6323 4156
rect 6349 4004 6355 4136
rect 6429 4104 6435 4236
rect 6445 4184 6451 4257
rect 6461 4144 6467 4196
rect 6493 4184 6499 4256
rect 6509 4224 6515 4256
rect 6525 4144 6531 4176
rect 6557 4144 6563 4216
rect 6573 4204 6579 4256
rect 6621 4244 6627 4256
rect 6653 4224 6659 4256
rect 6589 4164 6595 4196
rect 6653 4164 6659 4196
rect 6669 4164 6675 4236
rect 6509 4104 6515 4116
rect 6429 3984 6435 4096
rect 6621 4084 6627 4096
rect 6237 3904 6243 3916
rect 6093 3757 6124 3763
rect 5965 3684 5971 3716
rect 5917 3524 5923 3656
rect 5901 3464 5907 3496
rect 5933 3464 5939 3596
rect 5949 3504 5955 3676
rect 5965 3624 5971 3636
rect 5981 3604 5987 3736
rect 5997 3484 6003 3516
rect 6013 3504 6019 3756
rect 6029 3737 6060 3743
rect 6029 3724 6035 3737
rect 6093 3723 6099 3757
rect 6084 3717 6099 3723
rect 6045 3704 6051 3716
rect 6109 3704 6115 3716
rect 6029 3604 6035 3696
rect 6125 3684 6131 3696
rect 6045 3624 6051 3676
rect 6061 3464 6067 3516
rect 5940 3457 5955 3463
rect 5901 3424 5907 3456
rect 5885 3324 5891 3376
rect 5853 3124 5859 3176
rect 5405 3064 5411 3116
rect 5485 3064 5491 3116
rect 5885 3104 5891 3296
rect 5901 3184 5907 3336
rect 5917 3104 5923 3336
rect 5933 3264 5939 3316
rect 5949 3224 5955 3457
rect 6077 3364 6083 3636
rect 6125 3544 6131 3676
rect 6093 3504 6099 3536
rect 6109 3344 6115 3496
rect 6125 3444 6131 3476
rect 6029 3264 6035 3316
rect 6029 3244 6035 3256
rect 6109 3224 6115 3296
rect 5933 3104 5939 3136
rect 4797 2904 4803 2916
rect 5021 2903 5027 2936
rect 5149 2924 5155 2936
rect 5165 2924 5171 2936
rect 5069 2904 5075 2916
rect 5005 2897 5027 2903
rect 4808 2806 4814 2814
rect 4822 2806 4828 2814
rect 4836 2806 4842 2814
rect 4850 2806 4856 2814
rect 4797 2744 4803 2776
rect 4893 2724 4899 2736
rect 4669 2704 4675 2716
rect 4717 2704 4723 2716
rect 4637 2664 4643 2676
rect 4557 2644 4563 2656
rect 4605 2604 4611 2636
rect 4621 2584 4627 2636
rect 4397 2524 4403 2536
rect 4397 2344 4403 2476
rect 4429 2464 4435 2556
rect 4445 2544 4451 2556
rect 4333 2324 4339 2336
rect 4269 2302 4275 2316
rect 4397 2304 4403 2336
rect 4413 2304 4419 2316
rect 4125 2163 4131 2236
rect 4237 2184 4243 2276
rect 4381 2244 4387 2276
rect 4125 2157 4147 2163
rect 3981 2064 3987 2076
rect 3933 1904 3939 1996
rect 3933 1804 3939 1876
rect 3860 1757 3875 1763
rect 3677 1724 3683 1736
rect 3725 1723 3731 1736
rect 3757 1724 3763 1756
rect 3725 1717 3747 1723
rect 3581 1644 3587 1716
rect 3741 1703 3747 1717
rect 3741 1697 3756 1703
rect 3869 1664 3875 1757
rect 3901 1704 3907 1736
rect 3949 1664 3955 1736
rect 3597 1544 3603 1556
rect 3677 1504 3683 1616
rect 3476 1297 3491 1303
rect 2797 1124 2803 1196
rect 2829 1104 2835 1116
rect 2845 1064 2851 1236
rect 3149 1184 3155 1296
rect 3213 1243 3219 1296
rect 3197 1237 3219 1243
rect 3197 1184 3203 1237
rect 3277 1184 3283 1276
rect 3396 1237 3411 1243
rect 2877 1064 2883 1156
rect 3405 1144 3411 1237
rect 3437 1184 3443 1296
rect 3389 1104 3395 1116
rect 3213 1097 3228 1103
rect 2909 1064 2915 1076
rect 2717 1024 2723 1056
rect 2781 1044 2787 1056
rect 2717 964 2723 976
rect 2637 944 2643 956
rect 2580 897 2595 903
rect 2573 764 2579 896
rect 2621 844 2627 936
rect 2573 664 2579 736
rect 2605 724 2611 836
rect 2621 703 2627 836
rect 2637 784 2643 916
rect 2749 784 2755 896
rect 2685 704 2691 736
rect 2701 704 2707 716
rect 2621 697 2643 703
rect 2413 544 2419 576
rect 2477 564 2483 636
rect 2557 544 2563 656
rect 2013 443 2019 496
rect 2029 464 2035 516
rect 2333 504 2339 536
rect 2397 484 2403 516
rect 2013 437 2035 443
rect 1757 164 1763 276
rect 1805 184 1811 276
rect 1821 124 1827 296
rect 2029 283 2035 437
rect 2061 324 2067 436
rect 2477 343 2483 536
rect 2605 524 2611 696
rect 2621 604 2627 676
rect 2637 584 2643 697
rect 2749 684 2755 696
rect 2717 664 2723 676
rect 2669 584 2675 596
rect 2637 564 2643 576
rect 2749 564 2755 596
rect 2765 564 2771 596
rect 2509 504 2515 518
rect 2573 504 2579 516
rect 2685 504 2691 516
rect 2685 484 2691 496
rect 2461 337 2483 343
rect 2381 304 2387 316
rect 2413 304 2419 316
rect 2013 277 2035 283
rect 1869 224 1875 276
rect 1885 244 1891 276
rect 1853 124 1859 156
rect 1869 144 1875 216
rect 1885 124 1891 236
rect 1757 84 1763 96
rect 1869 84 1875 116
rect 1901 104 1907 176
rect 1933 104 1939 236
rect 1949 104 1955 236
rect 2013 184 2019 277
rect 1965 144 1971 156
rect 1997 144 2003 176
rect 2029 144 2035 176
rect 2077 144 2083 294
rect 2157 284 2163 296
rect 2317 204 2323 236
rect 2109 144 2115 176
rect 2237 164 2243 196
rect 2317 177 2332 183
rect 1981 104 1987 116
rect 2045 104 2051 116
rect 2125 104 2131 156
rect 2173 143 2179 156
rect 2173 137 2195 143
rect 2237 140 2243 156
rect 2317 144 2323 177
rect 2429 144 2435 256
rect 2461 164 2467 337
rect 2589 324 2595 356
rect 2477 264 2483 276
rect 2509 184 2515 276
rect 2557 263 2563 296
rect 2541 257 2563 263
rect 2541 184 2547 257
rect 2189 124 2195 137
rect 2253 104 2259 136
rect 2317 124 2323 136
rect 2461 104 2467 118
rect 2557 104 2563 176
rect 2573 164 2579 276
rect 2605 203 2611 316
rect 2669 304 2675 336
rect 2701 324 2707 436
rect 2701 284 2707 316
rect 2717 304 2723 556
rect 2797 524 2803 696
rect 2813 564 2819 1036
rect 2845 924 2851 1056
rect 2909 984 2915 1016
rect 2845 744 2851 916
rect 2829 704 2835 716
rect 2845 704 2851 716
rect 2861 697 2876 703
rect 2845 644 2851 656
rect 2861 584 2867 697
rect 2877 504 2883 596
rect 2893 584 2899 956
rect 2957 944 2963 1036
rect 3005 904 3011 936
rect 3053 924 3059 976
rect 3069 944 3075 956
rect 3069 864 3075 936
rect 2909 523 2915 856
rect 3053 744 3059 836
rect 3085 784 3091 1076
rect 3213 1064 3219 1097
rect 3117 904 3123 976
rect 3213 964 3219 1056
rect 3229 984 3235 1076
rect 3245 924 3251 1096
rect 3357 1044 3363 1076
rect 3341 1037 3356 1043
rect 3272 1006 3278 1014
rect 3286 1006 3292 1014
rect 3300 1006 3306 1014
rect 3314 1006 3320 1014
rect 3261 904 3267 936
rect 3181 824 3187 896
rect 3293 884 3299 916
rect 3341 904 3347 1037
rect 3389 883 3395 1096
rect 3485 1084 3491 1297
rect 3501 1284 3507 1336
rect 3501 1203 3507 1276
rect 3565 1204 3571 1476
rect 3597 1384 3603 1456
rect 3709 1443 3715 1596
rect 3725 1544 3731 1636
rect 3741 1544 3747 1656
rect 3933 1504 3939 1536
rect 3965 1504 3971 1636
rect 3981 1564 3987 2036
rect 3997 2023 4003 2096
rect 4061 2084 4067 2096
rect 3997 2017 4019 2023
rect 4013 1944 4019 2017
rect 3997 1724 4003 1816
rect 4013 1744 4019 1936
rect 4045 1924 4051 2036
rect 4061 1884 4067 2076
rect 4061 1804 4067 1856
rect 4077 1824 4083 1956
rect 4093 1924 4099 2116
rect 4141 1984 4147 2157
rect 4157 1884 4163 1996
rect 4173 1904 4179 2156
rect 4237 2144 4243 2176
rect 4333 2124 4339 2236
rect 4413 2224 4419 2276
rect 4189 1904 4195 1916
rect 4237 1904 4243 2056
rect 4061 1784 4067 1796
rect 4109 1744 4115 1876
rect 4221 1864 4227 1896
rect 4285 1884 4291 1976
rect 4317 1884 4323 1936
rect 4141 1744 4147 1836
rect 4269 1804 4275 1836
rect 4349 1784 4355 2216
rect 4429 2143 4435 2436
rect 4461 2304 4467 2576
rect 4541 2524 4547 2556
rect 4477 2504 4483 2516
rect 4477 2484 4483 2496
rect 4525 2484 4531 2516
rect 4541 2504 4547 2516
rect 4557 2504 4563 2556
rect 4445 2284 4451 2296
rect 4477 2264 4483 2476
rect 4509 2384 4515 2476
rect 4509 2344 4515 2376
rect 4525 2324 4531 2436
rect 4557 2344 4563 2476
rect 4589 2424 4595 2536
rect 4589 2344 4595 2396
rect 4461 2184 4467 2236
rect 4477 2204 4483 2256
rect 4493 2224 4499 2316
rect 4541 2264 4547 2276
rect 4445 2164 4451 2176
rect 4429 2137 4451 2143
rect 4413 1984 4419 2136
rect 4365 1864 4371 1916
rect 4445 1904 4451 2137
rect 4493 2124 4499 2176
rect 4509 1984 4515 2256
rect 4541 2223 4547 2256
rect 4557 2244 4563 2316
rect 4573 2304 4579 2316
rect 4605 2283 4611 2576
rect 4637 2544 4643 2556
rect 4653 2524 4659 2616
rect 4749 2526 4755 2536
rect 4669 2304 4675 2336
rect 4605 2277 4627 2283
rect 4621 2264 4627 2277
rect 4653 2264 4659 2276
rect 4685 2264 4691 2496
rect 4765 2484 4771 2636
rect 4829 2604 4835 2676
rect 4717 2284 4723 2396
rect 4765 2284 4771 2456
rect 4781 2343 4787 2596
rect 4808 2406 4814 2414
rect 4822 2406 4828 2414
rect 4836 2406 4842 2414
rect 4850 2406 4856 2414
rect 4781 2337 4803 2343
rect 4525 2217 4547 2223
rect 4525 2184 4531 2217
rect 4541 2164 4547 2196
rect 4557 2184 4563 2236
rect 4573 2224 4579 2236
rect 4653 2224 4659 2256
rect 4589 2184 4595 2196
rect 4573 1984 4579 2116
rect 4509 1904 4515 1916
rect 4397 1884 4403 1896
rect 4253 1726 4259 1776
rect 4381 1744 4387 1756
rect 4365 1724 4371 1736
rect 4013 1544 4019 1676
rect 4077 1644 4083 1716
rect 4189 1684 4195 1716
rect 4397 1704 4403 1796
rect 4413 1744 4419 1836
rect 4445 1743 4451 1796
rect 4461 1764 4467 1876
rect 4621 1864 4627 1896
rect 4637 1884 4643 2016
rect 4653 1884 4659 2216
rect 4717 2126 4723 2196
rect 4797 2184 4803 2337
rect 4813 2304 4819 2376
rect 4877 2364 4883 2436
rect 4829 2304 4835 2316
rect 4829 2284 4835 2296
rect 4845 2244 4851 2316
rect 4797 2164 4803 2176
rect 4781 1904 4787 2136
rect 4808 2006 4814 2014
rect 4822 2006 4828 2014
rect 4836 2006 4842 2014
rect 4850 2006 4856 2014
rect 4772 1877 4787 1883
rect 4477 1804 4483 1836
rect 4445 1737 4460 1743
rect 4493 1704 4499 1736
rect 4525 1726 4531 1836
rect 4541 1824 4547 1856
rect 4557 1844 4563 1856
rect 4077 1604 4083 1636
rect 4413 1604 4419 1696
rect 4557 1643 4563 1836
rect 4621 1724 4627 1856
rect 4637 1764 4643 1876
rect 4765 1844 4771 1856
rect 4781 1844 4787 1877
rect 4813 1864 4819 1896
rect 4877 1884 4883 1936
rect 4893 1904 4899 1936
rect 4653 1784 4659 1796
rect 4685 1784 4691 1816
rect 4541 1637 4563 1643
rect 4093 1583 4099 1596
rect 4084 1577 4099 1583
rect 4253 1544 4259 1556
rect 3700 1437 3715 1443
rect 3597 1364 3603 1376
rect 3501 1197 3523 1203
rect 3453 984 3459 1076
rect 3469 1044 3475 1056
rect 3380 877 3395 883
rect 3405 864 3411 936
rect 3501 924 3507 1096
rect 3517 984 3523 1197
rect 3549 1104 3555 1136
rect 3597 1084 3603 1176
rect 3565 984 3571 1036
rect 3613 944 3619 1056
rect 3629 984 3635 1116
rect 3693 1084 3699 1136
rect 3709 1104 3715 1437
rect 3741 1324 3747 1336
rect 3773 1163 3779 1476
rect 3853 1464 3859 1496
rect 3885 1464 3891 1476
rect 3789 1424 3795 1456
rect 3805 1404 3811 1436
rect 3837 1384 3843 1416
rect 3917 1384 3923 1476
rect 3981 1384 3987 1456
rect 4045 1384 4051 1516
rect 4061 1464 4067 1476
rect 4109 1464 4115 1476
rect 4077 1424 4083 1456
rect 4093 1384 4099 1416
rect 3821 1364 3827 1376
rect 3869 1324 3875 1356
rect 3789 1224 3795 1316
rect 3757 1157 3779 1163
rect 3693 1064 3699 1076
rect 3709 1044 3715 1076
rect 3437 884 3443 896
rect 3069 777 3084 783
rect 2941 704 2947 736
rect 3005 704 3011 736
rect 3037 684 3043 696
rect 3069 544 3075 777
rect 3133 684 3139 776
rect 3357 704 3363 836
rect 3373 724 3379 816
rect 3613 724 3619 936
rect 3645 864 3651 896
rect 3661 784 3667 916
rect 3380 717 3395 723
rect 3389 704 3395 717
rect 3341 684 3347 696
rect 3133 564 3139 656
rect 3197 564 3203 596
rect 2909 517 2924 523
rect 2813 364 2819 476
rect 2957 444 2963 496
rect 2813 324 2819 356
rect 2605 197 2620 203
rect 2605 104 2611 136
rect 2621 124 2627 196
rect 2637 164 2643 276
rect 2637 144 2643 156
rect 2733 144 2739 256
rect 2749 184 2755 296
rect 2781 283 2787 316
rect 2813 284 2819 296
rect 2829 284 2835 356
rect 2845 304 2851 376
rect 2861 324 2867 336
rect 2893 324 2899 416
rect 2957 384 2963 436
rect 2772 277 2787 283
rect 2765 264 2771 276
rect 2797 223 2803 236
rect 2797 217 2819 223
rect 2749 144 2755 176
rect 2781 124 2787 156
rect 2813 104 2819 217
rect 2829 184 2835 256
rect 2893 164 2899 316
rect 2909 304 2915 336
rect 2925 184 2931 336
rect 2957 304 2963 336
rect 2989 304 2995 436
rect 2989 264 2995 296
rect 3005 184 3011 296
rect 3053 284 3059 396
rect 3117 384 3123 436
rect 3069 264 3075 296
rect 3101 284 3107 376
rect 3181 324 3187 436
rect 3133 284 3139 294
rect 3165 244 3171 276
rect 2893 144 2899 156
rect 2845 124 2851 136
rect 2925 124 2931 176
rect 2845 104 2851 116
rect 2957 104 2963 176
rect 3165 164 3171 236
rect 3245 164 3251 636
rect 3272 606 3278 614
rect 3286 606 3292 614
rect 3300 606 3306 614
rect 3314 606 3320 614
rect 3517 544 3523 656
rect 3629 584 3635 716
rect 3645 604 3651 636
rect 3645 564 3651 576
rect 3261 384 3267 436
rect 3341 384 3347 516
rect 3341 304 3347 356
rect 3272 206 3278 214
rect 3286 206 3292 214
rect 3300 206 3306 214
rect 3314 206 3320 214
rect 3389 184 3395 236
rect 3021 144 3027 156
rect 3405 144 3411 276
rect 3437 263 3443 436
rect 3661 424 3667 636
rect 3677 383 3683 856
rect 3709 724 3715 936
rect 3709 664 3715 716
rect 3709 543 3715 636
rect 3725 584 3731 1076
rect 3741 984 3747 1016
rect 3741 684 3747 956
rect 3757 944 3763 1157
rect 3869 1084 3875 1316
rect 3885 1284 3891 1336
rect 3933 1284 3939 1356
rect 4077 1344 4083 1376
rect 4109 1344 4115 1416
rect 4125 1324 4131 1336
rect 3885 1164 3891 1276
rect 3981 1184 3987 1296
rect 4045 1284 4051 1296
rect 3885 1064 3891 1096
rect 3981 1084 3987 1096
rect 4013 1084 4019 1116
rect 3837 984 3843 1036
rect 3933 1004 3939 1076
rect 4029 1064 4035 1096
rect 4093 1084 4099 1156
rect 3805 944 3811 956
rect 3853 944 3859 956
rect 3933 904 3939 976
rect 3949 944 3955 976
rect 3965 924 3971 1016
rect 3757 684 3763 896
rect 3837 884 3843 896
rect 3837 784 3843 876
rect 3789 704 3795 756
rect 3885 704 3891 876
rect 3917 864 3923 896
rect 3741 584 3747 656
rect 3789 644 3795 696
rect 3901 684 3907 716
rect 3933 684 3939 696
rect 3965 664 3971 796
rect 3981 684 3987 976
rect 4077 943 4083 1056
rect 4125 964 4131 1316
rect 4157 1284 4163 1496
rect 4173 1484 4179 1516
rect 4365 1504 4371 1516
rect 4205 1484 4211 1496
rect 4301 1424 4307 1476
rect 4285 1417 4300 1423
rect 4189 1304 4195 1316
rect 4205 1304 4211 1396
rect 4189 1184 4195 1296
rect 4221 1284 4227 1316
rect 4269 1284 4275 1336
rect 4285 1324 4291 1417
rect 4349 1384 4355 1496
rect 4333 1324 4339 1336
rect 4349 1324 4355 1336
rect 4365 1324 4371 1476
rect 4381 1324 4387 1496
rect 4429 1464 4435 1516
rect 4445 1464 4451 1476
rect 4461 1424 4467 1436
rect 4429 1384 4435 1396
rect 4324 1297 4348 1303
rect 4237 1264 4243 1276
rect 4237 1184 4243 1216
rect 4141 944 4147 1056
rect 4068 937 4083 943
rect 3997 864 4003 896
rect 4029 704 4035 856
rect 4077 684 4083 937
rect 4157 924 4163 1076
rect 4189 1024 4195 1036
rect 4221 984 4227 1176
rect 4253 1104 4259 1236
rect 4237 1044 4243 1076
rect 4285 1043 4291 1096
rect 4285 1037 4307 1043
rect 4269 964 4275 1016
rect 4109 904 4115 916
rect 4141 903 4147 916
rect 4132 897 4147 903
rect 4109 824 4115 836
rect 4109 784 4115 796
rect 4141 724 4147 897
rect 4157 724 4163 916
rect 4205 884 4211 956
rect 4269 944 4275 956
rect 4301 944 4307 1037
rect 4317 944 4323 1276
rect 4381 1264 4387 1296
rect 4397 1243 4403 1336
rect 4461 1324 4467 1416
rect 4493 1404 4499 1496
rect 4493 1337 4508 1343
rect 4493 1264 4499 1337
rect 4525 1304 4531 1316
rect 4381 1237 4403 1243
rect 4381 984 4387 1237
rect 4493 1184 4499 1256
rect 4525 1104 4531 1136
rect 4461 984 4467 1036
rect 4477 1024 4483 1036
rect 4509 1024 4515 1056
rect 4380 950 4388 956
rect 4413 944 4419 976
rect 4429 944 4435 956
rect 4269 784 4275 916
rect 4301 904 4307 936
rect 4237 704 4243 736
rect 4269 724 4275 776
rect 4093 684 4099 696
rect 3693 537 3715 543
rect 3693 524 3699 537
rect 3757 404 3763 636
rect 3805 484 3811 516
rect 3853 504 3859 636
rect 3949 524 3955 636
rect 4029 544 4035 616
rect 4125 564 4131 576
rect 4221 544 4227 596
rect 4253 584 4259 656
rect 4269 584 4275 716
rect 4285 704 4291 836
rect 4301 804 4307 896
rect 4285 563 4291 656
rect 4276 557 4291 563
rect 4173 484 4179 516
rect 3661 377 3683 383
rect 3629 264 3635 296
rect 3645 284 3651 376
rect 3661 324 3667 377
rect 3677 264 3683 296
rect 3437 257 3452 263
rect 3693 243 3699 336
rect 3757 284 3763 376
rect 3773 304 3779 456
rect 3917 304 3923 336
rect 3773 264 3779 296
rect 3677 237 3699 243
rect 3421 164 3427 176
rect 3533 164 3539 236
rect 3677 184 3683 237
rect 3709 224 3715 256
rect 3709 184 3715 216
rect 3725 164 3731 176
rect 3133 124 3139 136
rect 3453 124 3459 136
rect 3533 126 3539 136
rect 3693 124 3699 156
rect 3741 144 3747 256
rect 3869 244 3875 296
rect 3885 264 3891 296
rect 3901 284 3907 296
rect 3917 264 3923 276
rect 3821 184 3827 236
rect 3821 124 3827 136
rect 3837 124 3843 216
rect 3853 144 3859 156
rect 3885 144 3891 256
rect 3917 124 3923 216
rect 3933 184 3939 256
rect 3949 164 3955 436
rect 4029 284 4035 356
rect 3981 264 3987 276
rect 3949 124 3955 156
rect 3469 104 3475 116
rect 1997 83 2003 96
rect 2061 84 2067 96
rect 3661 84 3667 116
rect 3821 104 3827 116
rect 3869 104 3875 116
rect 3997 104 4003 276
rect 4045 263 4051 296
rect 4125 284 4131 476
rect 4205 464 4211 496
rect 4253 304 4259 556
rect 4301 544 4307 676
rect 4317 664 4323 696
rect 4381 684 4387 916
rect 4461 904 4467 956
rect 4477 924 4483 976
rect 4509 924 4515 956
rect 4525 924 4531 1096
rect 4541 884 4547 1637
rect 4701 1544 4707 1756
rect 4717 1644 4723 1716
rect 4589 1504 4595 1516
rect 4717 1504 4723 1636
rect 4749 1524 4755 1676
rect 4781 1584 4787 1836
rect 4813 1744 4819 1856
rect 4829 1824 4835 1856
rect 4909 1744 4915 2896
rect 4957 2704 4963 2856
rect 5005 2724 5011 2897
rect 4957 2564 4963 2696
rect 5005 2524 5011 2556
rect 5021 2524 5027 2876
rect 5069 2764 5075 2896
rect 5197 2864 5203 3056
rect 5341 3024 5347 3056
rect 5421 3024 5427 3056
rect 5533 3044 5539 3096
rect 5565 3064 5571 3076
rect 5261 2964 5267 2976
rect 5309 2864 5315 2936
rect 5357 2924 5363 2936
rect 5085 2664 5091 2716
rect 4925 2264 4931 2296
rect 4941 2284 4947 2336
rect 5005 2304 5011 2376
rect 4989 2284 4995 2296
rect 4957 2244 4963 2256
rect 4973 2204 4979 2236
rect 5037 2144 5043 2516
rect 5053 2404 5059 2456
rect 5053 2284 5059 2396
rect 5101 2304 5107 2836
rect 5277 2824 5283 2836
rect 5245 2704 5251 2796
rect 5133 2684 5139 2696
rect 5181 2644 5187 2676
rect 5165 2584 5171 2616
rect 5181 2584 5187 2636
rect 5229 2584 5235 2676
rect 5261 2664 5267 2696
rect 5181 2544 5187 2576
rect 5133 2404 5139 2536
rect 5213 2524 5219 2536
rect 5277 2524 5283 2816
rect 5293 2704 5299 2796
rect 5309 2584 5315 2696
rect 5357 2684 5363 2736
rect 5389 2724 5395 2976
rect 5437 2924 5443 3036
rect 5485 2964 5491 2996
rect 5389 2684 5395 2716
rect 5437 2684 5443 2876
rect 5309 2504 5315 2576
rect 5405 2564 5411 2676
rect 5437 2664 5443 2676
rect 5357 2524 5363 2536
rect 5453 2524 5459 2836
rect 5485 2743 5491 2956
rect 5533 2944 5539 2956
rect 5501 2804 5507 2836
rect 5517 2824 5523 2916
rect 5517 2764 5523 2816
rect 5469 2737 5491 2743
rect 5469 2724 5475 2737
rect 5469 2704 5475 2716
rect 5517 2684 5523 2716
rect 5565 2704 5571 3036
rect 5597 3004 5603 3070
rect 5613 2964 5619 3036
rect 5661 2964 5667 2996
rect 5581 2904 5587 2916
rect 5581 2724 5587 2816
rect 5565 2684 5571 2696
rect 5581 2684 5587 2716
rect 5597 2704 5603 2796
rect 5485 2544 5491 2636
rect 5501 2524 5507 2536
rect 5405 2484 5411 2516
rect 5213 2384 5219 2396
rect 5085 2224 5091 2256
rect 5021 2084 5027 2096
rect 4957 1924 4963 2076
rect 5037 2063 5043 2116
rect 5085 2063 5091 2216
rect 5037 2057 5059 2063
rect 5053 1984 5059 2057
rect 5069 2057 5091 2063
rect 5069 1924 5075 2057
rect 5085 1924 5091 2036
rect 4957 1904 4963 1916
rect 5085 1904 5091 1916
rect 4829 1684 4835 1716
rect 4925 1684 4931 1836
rect 4989 1824 4995 1896
rect 5005 1884 5011 1896
rect 5005 1744 5011 1776
rect 4808 1606 4814 1614
rect 4822 1606 4828 1614
rect 4836 1606 4842 1614
rect 4850 1606 4856 1614
rect 4989 1584 4995 1676
rect 4893 1504 4899 1536
rect 4589 1104 4595 1496
rect 4765 1464 4771 1476
rect 4605 1324 4611 1416
rect 4669 1404 4675 1436
rect 4717 1344 4723 1376
rect 4605 1004 4611 1316
rect 4605 944 4611 956
rect 4557 904 4563 916
rect 4621 864 4627 1336
rect 4733 1324 4739 1396
rect 4749 1363 4755 1436
rect 4781 1384 4787 1436
rect 4813 1424 4819 1496
rect 4973 1464 4979 1476
rect 4973 1443 4979 1456
rect 4989 1444 4995 1456
rect 4973 1437 4988 1443
rect 4749 1357 4764 1363
rect 4781 1304 4787 1356
rect 4909 1344 4915 1356
rect 4877 1324 4883 1336
rect 4925 1324 4931 1436
rect 4957 1364 4963 1436
rect 5021 1424 5027 1776
rect 5037 1724 5043 1816
rect 5053 1804 5059 1896
rect 5037 1584 5043 1676
rect 5101 1484 5107 2136
rect 5117 2124 5123 2176
rect 5261 2124 5267 2196
rect 5149 1943 5155 2036
rect 5181 1984 5187 2076
rect 5309 2004 5315 2156
rect 5373 2124 5379 2236
rect 5389 2164 5395 2356
rect 5405 2304 5411 2476
rect 5453 2384 5459 2516
rect 5517 2364 5523 2536
rect 5405 2284 5411 2296
rect 5389 2144 5395 2156
rect 5437 2144 5443 2316
rect 5533 2284 5539 2676
rect 5549 2584 5555 2656
rect 5565 2544 5571 2596
rect 5565 2504 5571 2536
rect 5597 2304 5603 2676
rect 5613 2624 5619 2916
rect 5661 2884 5667 2956
rect 5677 2844 5683 3096
rect 5725 3044 5731 3056
rect 5645 2724 5651 2836
rect 5693 2764 5699 2876
rect 5709 2804 5715 2916
rect 5725 2904 5731 3036
rect 5757 2924 5763 2936
rect 5741 2904 5747 2916
rect 5725 2824 5731 2896
rect 5741 2744 5747 2876
rect 5757 2784 5763 2836
rect 5773 2704 5779 3036
rect 5805 3004 5811 3076
rect 5837 3044 5843 3056
rect 5837 3004 5843 3036
rect 5805 2984 5811 2996
rect 5821 2784 5827 2916
rect 5885 2724 5891 3096
rect 5917 2944 5923 3096
rect 5901 2924 5907 2936
rect 5853 2704 5859 2716
rect 5933 2704 5939 2736
rect 5693 2644 5699 2696
rect 5709 2684 5715 2696
rect 5821 2684 5827 2696
rect 5757 2664 5763 2676
rect 5709 2584 5715 2616
rect 5661 2564 5667 2576
rect 5725 2564 5731 2636
rect 5741 2564 5747 2656
rect 5773 2584 5779 2676
rect 5869 2664 5875 2696
rect 5949 2684 5955 2696
rect 5965 2684 5971 3216
rect 6125 3144 6131 3276
rect 6141 3124 6147 3796
rect 6173 3764 6179 3796
rect 6173 3504 6179 3576
rect 6189 3524 6195 3836
rect 6237 3624 6243 3756
rect 6269 3740 6275 3956
rect 6365 3864 6371 3876
rect 6253 3664 6259 3736
rect 6285 3684 6291 3856
rect 6344 3806 6350 3814
rect 6358 3806 6364 3814
rect 6372 3806 6378 3814
rect 6386 3806 6392 3814
rect 6493 3784 6499 3896
rect 6541 3864 6547 3956
rect 6413 3757 6483 3763
rect 6413 3744 6419 3757
rect 6477 3743 6483 3757
rect 6477 3737 6492 3743
rect 6301 3724 6307 3736
rect 6317 3704 6323 3736
rect 6445 3724 6451 3736
rect 6397 3663 6403 3696
rect 6260 3657 6275 3663
rect 6397 3657 6419 3663
rect 6189 3504 6195 3516
rect 6205 3484 6211 3536
rect 6237 3504 6243 3616
rect 6253 3504 6259 3556
rect 6269 3524 6275 3657
rect 6285 3584 6291 3596
rect 6269 3504 6275 3516
rect 6285 3504 6291 3556
rect 6301 3524 6307 3536
rect 6365 3484 6371 3496
rect 6157 3464 6163 3476
rect 6237 3464 6243 3476
rect 6157 3123 6163 3436
rect 6173 3204 6179 3236
rect 6157 3117 6172 3123
rect 5997 2984 6003 2996
rect 5661 2524 5667 2556
rect 5725 2544 5731 2556
rect 5757 2544 5763 2556
rect 5805 2524 5811 2636
rect 5917 2624 5923 2676
rect 5965 2544 5971 2676
rect 5981 2664 5987 2680
rect 6013 2664 6019 3036
rect 6109 2944 6115 3076
rect 6141 3044 6147 3056
rect 6189 2944 6195 3416
rect 6221 3403 6227 3436
rect 6344 3406 6350 3414
rect 6358 3406 6364 3414
rect 6372 3406 6378 3414
rect 6386 3406 6392 3414
rect 6205 3397 6227 3403
rect 6205 3104 6211 3397
rect 6333 3324 6339 3336
rect 6301 3304 6307 3318
rect 6237 3184 6243 3216
rect 6237 2984 6243 3116
rect 6269 3104 6275 3196
rect 6413 3164 6419 3657
rect 6461 3503 6467 3736
rect 6509 3724 6515 3736
rect 6493 3704 6499 3716
rect 6477 3504 6483 3516
rect 6452 3497 6467 3503
rect 6445 3464 6451 3496
rect 6477 3384 6483 3496
rect 6493 3464 6499 3696
rect 6525 3684 6531 3836
rect 6557 3784 6563 3916
rect 6621 3904 6627 3916
rect 6637 3824 6643 3836
rect 6573 3724 6579 3816
rect 6573 3684 6579 3716
rect 6589 3704 6595 3756
rect 6621 3664 6627 3716
rect 6653 3624 6659 4156
rect 6685 4124 6691 4156
rect 6701 4084 6707 4096
rect 6669 3944 6675 3996
rect 6733 3964 6739 4136
rect 6781 4104 6787 4216
rect 6813 4124 6819 4536
rect 6829 4324 6835 4536
rect 6861 4504 6867 4516
rect 6829 4284 6835 4316
rect 6845 4304 6851 4496
rect 6861 4324 6867 4336
rect 6877 4323 6883 4496
rect 6868 4317 6883 4323
rect 6845 4164 6851 4236
rect 6925 4224 6931 4276
rect 6845 4064 6851 4118
rect 6733 3904 6739 3956
rect 6829 3904 6835 4036
rect 6669 3784 6675 3896
rect 6717 3884 6723 3896
rect 6685 3784 6691 3796
rect 6861 3784 6867 3896
rect 6893 3884 6899 4116
rect 6941 4084 6947 4536
rect 6957 4264 6963 4336
rect 6957 4183 6963 4256
rect 6973 4204 6979 4236
rect 6957 4177 6972 4183
rect 6989 4163 6995 4236
rect 7053 4184 7059 4436
rect 7117 4344 7123 4516
rect 7133 4444 7139 4536
rect 7149 4444 7155 4656
rect 7197 4564 7203 4636
rect 7213 4624 7219 4656
rect 7165 4544 7171 4556
rect 7245 4544 7251 4676
rect 7437 4584 7443 4696
rect 7357 4564 7363 4576
rect 7197 4424 7203 4536
rect 7277 4504 7283 4556
rect 7117 4302 7123 4316
rect 7149 4284 7155 4416
rect 7261 4324 7267 4336
rect 7277 4324 7283 4496
rect 7197 4284 7203 4296
rect 6973 4157 6995 4163
rect 6973 4084 6979 4157
rect 7085 4144 7091 4216
rect 7117 4184 7123 4256
rect 7149 4244 7155 4276
rect 7213 4264 7219 4296
rect 7229 4284 7235 4316
rect 7229 4184 7235 4256
rect 7261 4224 7267 4276
rect 7101 4164 7107 4176
rect 7261 4164 7267 4216
rect 7293 4184 7299 4336
rect 7309 4184 7315 4276
rect 7101 4144 7107 4156
rect 7085 3904 7091 3916
rect 6909 3784 6915 3836
rect 6525 3544 6531 3576
rect 6509 3484 6515 3516
rect 6525 3464 6531 3496
rect 6525 3384 6531 3436
rect 6445 3344 6451 3376
rect 6493 3303 6499 3356
rect 6541 3344 6547 3476
rect 6573 3444 6579 3496
rect 6605 3484 6611 3496
rect 6701 3464 6707 3536
rect 6669 3384 6675 3416
rect 6653 3344 6659 3376
rect 6701 3364 6707 3456
rect 6733 3384 6739 3716
rect 6749 3423 6755 3456
rect 6749 3417 6771 3423
rect 6701 3340 6707 3356
rect 6765 3344 6771 3417
rect 6781 3384 6787 3736
rect 6941 3724 6947 3736
rect 6813 3704 6819 3716
rect 6829 3664 6835 3716
rect 6829 3584 6835 3656
rect 6829 3504 6835 3576
rect 6861 3544 6867 3716
rect 6893 3704 6899 3716
rect 6909 3564 6915 3676
rect 6493 3297 6508 3303
rect 6509 3204 6515 3296
rect 6557 3224 6563 3336
rect 6765 3324 6771 3336
rect 6397 3104 6403 3116
rect 6205 2763 6211 2916
rect 6253 2904 6259 2916
rect 6189 2757 6211 2763
rect 6045 2584 6051 2696
rect 6093 2684 6099 2696
rect 6141 2664 6147 2696
rect 6164 2677 6179 2683
rect 5949 2537 5964 2543
rect 5613 2504 5619 2516
rect 5933 2504 5939 2516
rect 5949 2504 5955 2537
rect 5981 2504 5987 2516
rect 6013 2504 6019 2556
rect 6029 2504 6035 2516
rect 6061 2504 6067 2596
rect 6125 2544 6131 2576
rect 6141 2564 6147 2636
rect 6173 2524 6179 2677
rect 6173 2504 6179 2516
rect 5885 2464 5891 2496
rect 5917 2464 5923 2476
rect 5597 2284 5603 2296
rect 5485 2204 5491 2276
rect 5533 2264 5539 2276
rect 5341 2097 5356 2103
rect 5133 1937 5155 1943
rect 5133 1904 5139 1937
rect 5117 1804 5123 1896
rect 5133 1884 5139 1896
rect 5197 1844 5203 1876
rect 5229 1864 5235 1896
rect 5277 1884 5283 1896
rect 5245 1844 5251 1856
rect 5220 1837 5235 1843
rect 5117 1502 5123 1516
rect 5053 1344 5059 1476
rect 4749 1164 4755 1236
rect 4653 1102 4659 1116
rect 4740 1097 4755 1103
rect 4685 924 4691 936
rect 4701 924 4707 996
rect 4733 984 4739 1056
rect 4749 1044 4755 1097
rect 4765 1084 4771 1096
rect 4653 864 4659 896
rect 4413 702 4419 816
rect 4541 784 4547 796
rect 4685 684 4691 694
rect 4349 564 4355 636
rect 4381 624 4387 676
rect 4029 257 4051 263
rect 4013 164 4019 236
rect 4029 184 4035 257
rect 4173 164 4179 276
rect 4301 264 4307 296
rect 4317 284 4323 556
rect 4397 524 4403 536
rect 4045 124 4051 136
rect 4061 104 4067 156
rect 4109 144 4115 156
rect 4173 126 4179 136
rect 4093 104 4099 116
rect 4285 104 4291 236
rect 4333 223 4339 496
rect 4349 384 4355 456
rect 4420 437 4435 443
rect 4429 344 4435 437
rect 4429 324 4435 336
rect 4365 304 4371 316
rect 4445 304 4451 496
rect 4509 384 4515 476
rect 4461 304 4467 316
rect 4557 304 4563 436
rect 4429 283 4435 296
rect 4429 277 4451 283
rect 4333 217 4348 223
rect 4301 184 4307 196
rect 4333 164 4339 196
rect 4349 144 4355 216
rect 4365 184 4371 256
rect 4381 144 4387 256
rect 4445 184 4451 277
rect 4461 183 4467 296
rect 4525 277 4540 283
rect 4493 264 4499 276
rect 4509 243 4515 276
rect 4525 264 4531 277
rect 4493 237 4515 243
rect 4493 184 4499 237
rect 4525 184 4531 256
rect 4461 177 4483 183
rect 4461 104 4467 156
rect 4477 104 4483 177
rect 4557 164 4563 296
rect 4573 264 4579 336
rect 4621 324 4627 336
rect 4637 324 4643 356
rect 4653 324 4659 676
rect 4685 544 4691 656
rect 4669 464 4675 516
rect 4701 384 4707 616
rect 4765 524 4771 996
rect 4781 964 4787 1296
rect 4861 1264 4867 1316
rect 4941 1284 4947 1336
rect 5149 1323 5155 1736
rect 5213 1704 5219 1816
rect 5229 1764 5235 1837
rect 5229 1704 5235 1756
rect 5245 1743 5251 1836
rect 5261 1804 5267 1836
rect 5261 1763 5267 1796
rect 5261 1757 5283 1763
rect 5245 1737 5260 1743
rect 5261 1724 5267 1736
rect 5277 1724 5283 1757
rect 5293 1744 5299 1836
rect 5309 1744 5315 1996
rect 5341 1884 5347 2097
rect 5437 2044 5443 2136
rect 5517 2124 5523 2176
rect 5549 2144 5555 2236
rect 5597 2184 5603 2256
rect 5613 2184 5619 2316
rect 5629 2304 5635 2316
rect 5645 2304 5651 2336
rect 5741 2304 5747 2356
rect 5757 2304 5763 2376
rect 5629 2184 5635 2276
rect 5645 2264 5651 2296
rect 5661 2264 5667 2276
rect 5661 2184 5667 2256
rect 5581 2044 5587 2156
rect 5645 2144 5651 2156
rect 5661 2104 5667 2176
rect 5677 2124 5683 2296
rect 5725 2264 5731 2276
rect 5741 2264 5747 2296
rect 5789 2164 5795 2276
rect 5693 2144 5699 2156
rect 5789 2084 5795 2136
rect 5805 2124 5811 2336
rect 5837 2304 5843 2356
rect 5853 2284 5859 2316
rect 5933 2304 5939 2436
rect 5869 2257 5884 2263
rect 5869 2144 5875 2257
rect 5885 2184 5891 2216
rect 5821 2124 5827 2136
rect 5869 2084 5875 2136
rect 5901 2104 5907 2236
rect 5917 2184 5923 2256
rect 5501 1924 5507 2036
rect 5389 1904 5395 1916
rect 5341 1824 5347 1856
rect 5357 1804 5363 1876
rect 5325 1764 5331 1796
rect 5325 1744 5331 1756
rect 5373 1744 5379 1856
rect 5405 1784 5411 1916
rect 5421 1884 5427 1896
rect 5453 1824 5459 1916
rect 5549 1864 5555 1896
rect 5725 1864 5731 1936
rect 5469 1804 5475 1836
rect 5341 1724 5347 1736
rect 5405 1684 5411 1718
rect 5261 1524 5267 1576
rect 5293 1504 5299 1636
rect 5405 1502 5411 1556
rect 5341 1484 5347 1496
rect 5437 1484 5443 1736
rect 5341 1424 5347 1456
rect 5197 1344 5203 1356
rect 5245 1324 5251 1356
rect 5309 1344 5315 1356
rect 5437 1344 5443 1396
rect 5453 1344 5459 1376
rect 5469 1344 5475 1476
rect 5485 1444 5491 1496
rect 5485 1384 5491 1436
rect 5501 1344 5507 1416
rect 5517 1344 5523 1856
rect 5533 1784 5539 1816
rect 5613 1804 5619 1836
rect 5629 1744 5635 1756
rect 5661 1744 5667 1796
rect 5604 1737 5619 1743
rect 5613 1723 5619 1737
rect 5709 1724 5715 1776
rect 5725 1724 5731 1836
rect 5757 1764 5763 1996
rect 5837 1904 5843 1916
rect 5853 1904 5859 2036
rect 5917 1984 5923 2036
rect 5949 1964 5955 2396
rect 6109 2364 6115 2436
rect 5885 1764 5891 1876
rect 5981 1844 5987 2356
rect 6189 2344 6195 2757
rect 6205 2624 6211 2736
rect 6237 2624 6243 2836
rect 6269 2744 6275 3076
rect 6285 2644 6291 3076
rect 6301 2784 6307 3076
rect 6317 2984 6323 3096
rect 6397 3064 6403 3096
rect 6429 3084 6435 3096
rect 6445 3084 6451 3156
rect 6717 3144 6723 3316
rect 6749 3164 6755 3176
rect 6461 3104 6467 3116
rect 6509 3104 6515 3136
rect 6669 3104 6675 3116
rect 6717 3104 6723 3136
rect 6724 3097 6732 3103
rect 6493 3083 6499 3096
rect 6493 3077 6508 3083
rect 6344 3006 6350 3014
rect 6358 3006 6364 3014
rect 6372 3006 6378 3014
rect 6386 3006 6392 3014
rect 6541 2964 6547 2976
rect 6509 2884 6515 2936
rect 6557 2903 6563 3036
rect 6573 2964 6579 3096
rect 6589 3064 6595 3096
rect 6749 3084 6755 3156
rect 6685 3024 6691 3076
rect 6717 3044 6723 3076
rect 6765 3063 6771 3316
rect 6781 3104 6787 3116
rect 6797 3064 6803 3436
rect 6813 3424 6819 3456
rect 6861 3324 6867 3536
rect 6957 3524 6963 3636
rect 6900 3517 6915 3523
rect 6909 3484 6915 3517
rect 6957 3504 6963 3516
rect 6877 3184 6883 3416
rect 6909 3384 6915 3476
rect 6973 3444 6979 3836
rect 6989 3684 6995 3696
rect 7021 3504 7027 3736
rect 7085 3484 7091 3496
rect 7021 3424 7027 3476
rect 6909 3344 6915 3376
rect 7021 3344 7027 3416
rect 7053 3384 7059 3456
rect 7069 3424 7075 3476
rect 7101 3404 7107 4116
rect 7165 4084 7171 4156
rect 7197 4124 7203 4136
rect 7181 4104 7187 4116
rect 7181 3784 7187 4016
rect 7261 3864 7267 4156
rect 7325 4144 7331 4296
rect 7373 4284 7379 4296
rect 7373 4224 7379 4276
rect 7389 4244 7395 4296
rect 7373 4144 7379 4196
rect 7389 4144 7395 4156
rect 7405 4143 7411 4556
rect 7421 4344 7427 4536
rect 7437 4364 7443 4496
rect 7453 4404 7459 5297
rect 7485 5164 7491 5356
rect 7517 5344 7523 5476
rect 7485 5044 7491 5156
rect 7501 5104 7507 5116
rect 7517 5084 7523 5336
rect 7565 5264 7571 5316
rect 7485 4704 7491 4716
rect 7485 4544 7491 4556
rect 7437 4264 7443 4316
rect 7453 4284 7459 4296
rect 7469 4284 7475 4536
rect 7501 4524 7507 5076
rect 7517 4944 7523 5076
rect 7517 4704 7523 4756
rect 7533 4684 7539 4736
rect 7565 4624 7571 4636
rect 7581 4604 7587 5718
rect 7693 5504 7699 5736
rect 7709 5644 7715 5716
rect 7757 5502 7763 5536
rect 7693 5484 7699 5496
rect 7821 5484 7827 5636
rect 7837 5624 7843 5736
rect 7869 5544 7875 5556
rect 7885 5544 7891 5556
rect 7917 5524 7923 5536
rect 7613 5424 7619 5456
rect 7693 5324 7699 5436
rect 7780 5337 7795 5343
rect 7629 5064 7635 5136
rect 7693 5084 7699 5316
rect 7741 5304 7747 5336
rect 7789 5304 7795 5337
rect 7821 5304 7827 5456
rect 7837 5444 7843 5456
rect 7837 5344 7843 5436
rect 7901 5384 7907 5496
rect 7949 5464 7955 5496
rect 7949 5324 7955 5416
rect 7965 5364 7971 5476
rect 7709 5124 7715 5136
rect 7741 5104 7747 5236
rect 7773 5184 7779 5256
rect 7629 5024 7635 5056
rect 7725 5024 7731 5056
rect 7613 4904 7619 4996
rect 7741 4964 7747 5056
rect 7773 5004 7779 5096
rect 7789 4964 7795 5296
rect 7805 5284 7811 5296
rect 7853 5284 7859 5316
rect 7821 5244 7827 5276
rect 7853 5164 7859 5236
rect 7805 5124 7811 5156
rect 7853 5104 7859 5116
rect 7869 5104 7875 5236
rect 7901 5124 7907 5316
rect 7933 5104 7939 5116
rect 7821 5064 7827 5076
rect 7613 4884 7619 4896
rect 7629 4844 7635 4916
rect 7645 4884 7651 4896
rect 7597 4684 7603 4776
rect 7677 4744 7683 4916
rect 7725 4904 7731 4916
rect 7693 4784 7699 4836
rect 7709 4744 7715 4756
rect 7636 4697 7651 4703
rect 7549 4544 7555 4556
rect 7645 4544 7651 4697
rect 7677 4544 7683 4656
rect 7725 4644 7731 4856
rect 7741 4704 7747 4956
rect 7821 4944 7827 5036
rect 7741 4664 7747 4696
rect 7757 4684 7763 4736
rect 7805 4704 7811 4916
rect 7821 4724 7827 4936
rect 7837 4884 7843 4896
rect 7853 4783 7859 5076
rect 7917 4984 7923 5076
rect 7933 4964 7939 5076
rect 7949 5004 7955 5096
rect 7869 4937 7884 4943
rect 7869 4904 7875 4937
rect 7885 4897 7900 4903
rect 7869 4804 7875 4836
rect 7853 4777 7875 4783
rect 7853 4724 7859 4756
rect 7821 4684 7827 4716
rect 7853 4704 7859 4716
rect 7789 4664 7795 4676
rect 7533 4524 7539 4536
rect 7581 4504 7587 4536
rect 7645 4504 7651 4516
rect 7693 4504 7699 4616
rect 7773 4564 7779 4636
rect 7725 4524 7731 4556
rect 7741 4503 7747 4536
rect 7725 4497 7747 4503
rect 7396 4137 7411 4143
rect 7309 4104 7315 4116
rect 7309 3984 7315 4096
rect 7293 3884 7299 3936
rect 7357 3924 7363 4036
rect 7389 3923 7395 4136
rect 7437 4104 7443 4156
rect 7453 4084 7459 4256
rect 7469 4164 7475 4276
rect 7485 4164 7491 4436
rect 7501 4324 7507 4336
rect 7501 4244 7507 4296
rect 7469 4084 7475 4136
rect 7380 3917 7395 3923
rect 7373 3884 7379 3896
rect 7533 3884 7539 4416
rect 7581 4404 7587 4496
rect 7565 4284 7571 4356
rect 7565 4204 7571 4276
rect 7581 4264 7587 4296
rect 7549 4164 7555 4196
rect 7645 4164 7651 4496
rect 7693 4324 7699 4336
rect 7613 4104 7619 4116
rect 7661 4104 7667 4116
rect 7565 3904 7571 4036
rect 7613 3964 7619 4036
rect 7613 3924 7619 3956
rect 7309 3863 7315 3876
rect 7293 3857 7315 3863
rect 7181 3764 7187 3776
rect 7117 3684 7123 3718
rect 7149 3704 7155 3736
rect 7165 3584 7171 3676
rect 7181 3544 7187 3556
rect 7165 3484 7171 3496
rect 7133 3384 7139 3436
rect 7037 3344 7043 3376
rect 7069 3364 7075 3376
rect 7149 3364 7155 3396
rect 7197 3384 7203 3856
rect 7293 3703 7299 3857
rect 7309 3726 7315 3736
rect 7341 3704 7347 3736
rect 7293 3697 7315 3703
rect 7213 3464 7219 3616
rect 7309 3584 7315 3697
rect 7245 3524 7251 3536
rect 7213 3364 7219 3456
rect 7277 3404 7283 3456
rect 7277 3364 7283 3396
rect 6845 3104 6851 3136
rect 6877 3124 6883 3176
rect 6861 3104 6867 3116
rect 6749 3057 6771 3063
rect 6637 2964 6643 2976
rect 6573 2924 6579 2936
rect 6701 2924 6707 3036
rect 6557 2897 6572 2903
rect 6205 2544 6211 2576
rect 6237 2564 6243 2596
rect 6237 2544 6243 2556
rect 6253 2544 6259 2556
rect 6301 2524 6307 2696
rect 6333 2684 6339 2876
rect 6669 2783 6675 2876
rect 6669 2777 6691 2783
rect 6685 2684 6691 2777
rect 6733 2704 6739 2996
rect 6749 2944 6755 3057
rect 6765 3024 6771 3036
rect 6813 2983 6819 3036
rect 6845 3004 6851 3096
rect 6877 3024 6883 3116
rect 6813 2977 6835 2983
rect 6829 2944 6835 2977
rect 6893 2983 6899 3336
rect 7165 3284 7171 3316
rect 7293 3264 7299 3456
rect 7117 3204 7123 3236
rect 6909 3104 6915 3116
rect 6973 3104 6979 3156
rect 7037 3144 7043 3156
rect 7085 3124 7091 3196
rect 6989 3064 6995 3096
rect 6893 2977 6915 2983
rect 6845 2924 6851 2976
rect 6909 2964 6915 2977
rect 6893 2904 6899 2956
rect 6781 2684 6787 2696
rect 6909 2684 6915 2956
rect 6925 2924 6931 2996
rect 6941 2944 6947 3056
rect 6989 3037 6995 3056
rect 6941 2704 6947 2896
rect 6957 2784 6963 2896
rect 6973 2784 6979 2996
rect 6989 2944 6995 3016
rect 7037 2964 7043 3016
rect 7117 2964 7123 3116
rect 7133 3084 7139 3096
rect 7149 3044 7155 3116
rect 7005 2783 7011 2956
rect 7133 2944 7139 3016
rect 7229 2944 7235 3076
rect 7261 2984 7267 3096
rect 7341 3064 7347 3096
rect 7357 3084 7363 3316
rect 7357 2944 7363 3076
rect 7373 2944 7379 2956
rect 7389 2944 7395 3876
rect 7405 3864 7411 3876
rect 7421 3684 7427 3716
rect 7453 3704 7459 3736
rect 7469 3724 7475 3736
rect 7485 3704 7491 3876
rect 7533 3744 7539 3756
rect 7485 3504 7491 3696
rect 7565 3524 7571 3896
rect 7597 3744 7603 3756
rect 7581 3664 7587 3716
rect 7613 3704 7619 3836
rect 7645 3744 7651 3876
rect 7661 3764 7667 3836
rect 7677 3744 7683 3916
rect 7693 3904 7699 4236
rect 7709 3924 7715 4136
rect 7725 3943 7731 4497
rect 7789 4484 7795 4636
rect 7837 4524 7843 4656
rect 7853 4524 7859 4536
rect 7764 4437 7779 4443
rect 7773 4344 7779 4437
rect 7757 4323 7763 4336
rect 7757 4317 7795 4323
rect 7789 4304 7795 4317
rect 7773 4284 7779 4296
rect 7789 4144 7795 4216
rect 7773 4044 7779 4136
rect 7789 4084 7795 4116
rect 7805 4064 7811 4336
rect 7821 4304 7827 4316
rect 7837 4284 7843 4296
rect 7821 4024 7827 4276
rect 7837 4164 7843 4276
rect 7869 4243 7875 4777
rect 7885 4744 7891 4897
rect 7965 4884 7971 5356
rect 7981 5344 7987 5476
rect 7997 5424 8003 5496
rect 8013 5384 8019 5636
rect 8109 5484 8115 5496
rect 8125 5484 8131 5496
rect 8045 5444 8051 5456
rect 8077 5384 8083 5436
rect 8029 5364 8035 5376
rect 8141 5344 8147 5356
rect 7997 5324 8003 5336
rect 7981 5284 7987 5316
rect 8029 5304 8035 5336
rect 8013 5184 8019 5276
rect 7997 5064 8003 5116
rect 8061 5103 8067 5116
rect 8061 5097 8083 5103
rect 7997 5044 8003 5056
rect 7981 4940 7987 5016
rect 7997 4944 8003 4956
rect 8013 4944 8019 5056
rect 7901 4624 7907 4856
rect 7917 4664 7923 4676
rect 7965 4664 7971 4796
rect 7981 4663 7987 4932
rect 8045 4884 8051 4896
rect 8061 4744 8067 5076
rect 8077 4984 8083 5097
rect 8093 5084 8099 5096
rect 8093 4764 8099 4876
rect 8109 4864 8115 4956
rect 8125 4924 8131 5096
rect 7997 4684 8003 4716
rect 8125 4684 8131 4876
rect 8029 4664 8035 4676
rect 7981 4657 8003 4663
rect 7949 4584 7955 4656
rect 7901 4302 7907 4356
rect 7917 4284 7923 4536
rect 7981 4524 7987 4636
rect 7997 4604 8003 4657
rect 8013 4524 8019 4536
rect 7853 4237 7875 4243
rect 7837 4044 7843 4096
rect 7725 3937 7747 3943
rect 7693 3764 7699 3896
rect 7709 3884 7715 3896
rect 7700 3717 7724 3723
rect 7629 3704 7635 3716
rect 7645 3704 7651 3716
rect 7437 3464 7443 3496
rect 7485 3484 7491 3496
rect 7597 3364 7603 3516
rect 7693 3464 7699 3476
rect 7501 3344 7507 3356
rect 7613 3337 7644 3343
rect 7421 3284 7427 3318
rect 7485 3184 7491 3236
rect 7501 3184 7507 3316
rect 7517 3304 7523 3336
rect 7613 3324 7619 3337
rect 7661 3323 7667 3456
rect 7677 3404 7683 3436
rect 7645 3317 7667 3323
rect 7549 3284 7555 3316
rect 7533 3264 7539 3276
rect 7453 3124 7459 3156
rect 7485 3144 7491 3156
rect 7613 3124 7619 3296
rect 7629 3264 7635 3316
rect 7501 3104 7507 3116
rect 7421 3004 7427 3076
rect 7517 3004 7523 3116
rect 7533 3104 7539 3116
rect 7613 3104 7619 3116
rect 7629 3104 7635 3256
rect 7581 3084 7587 3096
rect 7597 3084 7603 3096
rect 7645 3084 7651 3317
rect 7661 3284 7667 3296
rect 7549 3064 7555 3076
rect 7645 3064 7651 3076
rect 7677 3064 7683 3336
rect 7693 3304 7699 3316
rect 7709 3303 7715 3396
rect 7725 3364 7731 3516
rect 7741 3363 7747 3937
rect 7757 3844 7763 3856
rect 7757 3724 7763 3836
rect 7773 3524 7779 3736
rect 7789 3724 7795 3956
rect 7821 3743 7827 4016
rect 7805 3737 7827 3743
rect 7789 3664 7795 3676
rect 7789 3584 7795 3656
rect 7805 3504 7811 3737
rect 7837 3724 7843 3736
rect 7853 3664 7859 4237
rect 7869 4064 7875 4076
rect 7885 4004 7891 4116
rect 7901 4104 7907 4116
rect 7901 4064 7907 4076
rect 7869 3744 7875 3756
rect 7885 3743 7891 3976
rect 7917 3884 7923 4276
rect 7933 3944 7939 4476
rect 7949 4404 7955 4436
rect 8029 4384 8035 4596
rect 8045 4384 8051 4616
rect 7949 4124 7955 4176
rect 7965 4084 7971 4136
rect 7949 3924 7955 4036
rect 7917 3744 7923 3876
rect 7965 3803 7971 4056
rect 7981 3964 7987 4096
rect 7997 3984 8003 4036
rect 7997 3904 8003 3956
rect 8013 3924 8019 4076
rect 7965 3797 7987 3803
rect 7885 3737 7900 3743
rect 7773 3484 7779 3496
rect 7757 3384 7763 3436
rect 7741 3357 7763 3363
rect 7741 3304 7747 3316
rect 7757 3304 7763 3357
rect 7773 3323 7779 3476
rect 7789 3344 7795 3396
rect 7773 3317 7795 3323
rect 7709 3297 7724 3303
rect 7789 3224 7795 3317
rect 7805 3264 7811 3296
rect 7821 3284 7827 3656
rect 7901 3504 7907 3516
rect 7949 3484 7955 3736
rect 7981 3726 7987 3797
rect 7981 3384 7987 3436
rect 7837 3344 7843 3356
rect 7949 3344 7955 3356
rect 7965 3304 7971 3356
rect 7997 3324 8003 3336
rect 7812 3257 7827 3263
rect 7725 3124 7731 3216
rect 7805 3104 7811 3116
rect 7821 3084 7827 3257
rect 7837 3104 7843 3156
rect 7764 3077 7779 3083
rect 7677 3004 7683 3056
rect 7709 2984 7715 3036
rect 7437 2944 7443 2956
rect 7085 2924 7091 2936
rect 6996 2777 7011 2783
rect 7117 2702 7123 2836
rect 7149 2724 7155 2816
rect 6344 2606 6350 2614
rect 6358 2606 6364 2614
rect 6372 2606 6378 2614
rect 6386 2606 6392 2614
rect 6413 2584 6419 2676
rect 6429 2584 6435 2636
rect 6445 2564 6451 2636
rect 6349 2544 6355 2556
rect 6525 2544 6531 2636
rect 6653 2584 6659 2676
rect 6749 2564 6755 2616
rect 6765 2604 6771 2636
rect 6781 2544 6787 2676
rect 6269 2504 6275 2516
rect 6308 2497 6323 2503
rect 6301 2384 6307 2476
rect 6285 2344 6291 2356
rect 6100 2337 6115 2343
rect 6109 2303 6115 2337
rect 6125 2324 6131 2336
rect 6317 2324 6323 2497
rect 6541 2484 6547 2516
rect 6589 2304 6595 2536
rect 6669 2484 6675 2496
rect 6109 2297 6124 2303
rect 6013 2224 6019 2296
rect 6077 2284 6083 2296
rect 6029 2164 6035 2276
rect 6077 2164 6083 2236
rect 6045 2126 6051 2156
rect 6109 2144 6115 2276
rect 6157 2244 6163 2296
rect 6189 2224 6195 2256
rect 6205 2144 6211 2276
rect 6461 2264 6467 2276
rect 6237 2140 6243 2156
rect 6109 2084 6115 2136
rect 6253 2024 6259 2256
rect 6344 2206 6350 2214
rect 6358 2206 6364 2214
rect 6372 2206 6378 2214
rect 6386 2206 6392 2214
rect 6333 2144 6339 2176
rect 6365 2144 6371 2156
rect 6413 2144 6419 2236
rect 6445 2224 6451 2256
rect 6541 2244 6547 2294
rect 6477 2164 6483 2236
rect 6525 2184 6531 2196
rect 6605 2184 6611 2476
rect 6653 2244 6659 2436
rect 6701 2384 6707 2516
rect 6445 2124 6451 2136
rect 6477 2123 6483 2156
rect 6541 2124 6547 2156
rect 6468 2117 6483 2123
rect 6317 2104 6323 2116
rect 6445 2084 6451 2096
rect 6477 2064 6483 2096
rect 5965 1764 5971 1796
rect 6013 1764 6019 1876
rect 5613 1717 5628 1723
rect 5597 1704 5603 1716
rect 5693 1584 5699 1636
rect 5933 1584 5939 1756
rect 6077 1724 6083 1956
rect 5981 1544 5987 1636
rect 5732 1537 5779 1543
rect 5693 1524 5699 1536
rect 5597 1517 5612 1523
rect 5597 1484 5603 1517
rect 5773 1504 5779 1537
rect 5805 1537 5875 1543
rect 5805 1504 5811 1537
rect 5828 1517 5852 1523
rect 5869 1504 5875 1537
rect 5693 1497 5708 1503
rect 5629 1484 5635 1496
rect 5133 1317 5155 1323
rect 4808 1206 4814 1214
rect 4822 1206 4828 1214
rect 4836 1206 4842 1214
rect 4850 1206 4856 1214
rect 4797 1084 4803 1156
rect 4797 1064 4803 1076
rect 4781 904 4787 916
rect 4797 864 4803 956
rect 4813 944 4819 1036
rect 4877 984 4883 1276
rect 4909 1104 4915 1116
rect 4909 1064 4915 1076
rect 4845 844 4851 876
rect 4861 844 4867 936
rect 4893 864 4899 936
rect 4909 924 4915 976
rect 4925 944 4931 1096
rect 4941 1024 4947 1236
rect 4989 1124 4995 1256
rect 5069 1184 5075 1196
rect 5053 1124 5059 1136
rect 5069 1084 5075 1096
rect 4996 1077 5011 1083
rect 4989 964 4995 1056
rect 5005 1004 5011 1077
rect 5021 1064 5027 1076
rect 5005 984 5011 996
rect 5021 964 5027 1016
rect 5069 984 5075 1076
rect 5085 1064 5091 1116
rect 5117 1084 5123 1096
rect 5101 1064 5107 1076
rect 5085 944 5091 1056
rect 4973 924 4979 936
rect 5101 924 5107 1016
rect 5133 904 5139 1317
rect 5149 1244 5155 1296
rect 5149 1224 5155 1236
rect 5165 1184 5171 1236
rect 5213 1184 5219 1276
rect 5325 1244 5331 1336
rect 5437 1264 5443 1316
rect 5277 1117 5292 1123
rect 5149 964 5155 996
rect 5165 984 5171 1116
rect 5261 1104 5267 1116
rect 5181 1064 5187 1096
rect 5181 1044 5187 1056
rect 5229 984 5235 1016
rect 5261 1004 5267 1096
rect 5277 1084 5283 1117
rect 5213 964 5219 976
rect 5293 964 5299 1076
rect 4781 704 4787 836
rect 4808 806 4814 814
rect 4822 806 4828 814
rect 4836 806 4842 814
rect 4850 806 4856 814
rect 4877 664 4883 676
rect 4909 584 4915 616
rect 4781 564 4787 576
rect 4957 564 4963 896
rect 5213 884 5219 956
rect 4989 784 4995 836
rect 5021 684 5027 876
rect 5133 764 5139 836
rect 5181 704 5187 716
rect 4989 564 4995 676
rect 5005 644 5011 656
rect 5037 584 5043 696
rect 5069 684 5075 696
rect 5085 624 5091 676
rect 5101 603 5107 696
rect 5197 684 5203 756
rect 5220 697 5235 703
rect 5085 597 5107 603
rect 4893 544 4899 556
rect 4808 406 4814 414
rect 4822 406 4828 414
rect 4836 406 4842 414
rect 4850 406 4856 414
rect 4941 364 4947 436
rect 4573 224 4579 256
rect 4509 144 4515 156
rect 4557 144 4563 156
rect 4589 144 4595 156
rect 4605 124 4611 296
rect 4621 224 4627 316
rect 4653 304 4659 316
rect 4685 264 4691 336
rect 4701 304 4707 316
rect 4653 184 4659 256
rect 4717 184 4723 316
rect 4733 284 4739 296
rect 4637 104 4643 136
rect 4685 124 4691 176
rect 4733 164 4739 276
rect 4701 104 4707 136
rect 4749 104 4755 136
rect 4813 104 4819 176
rect 4829 104 4835 276
rect 4861 144 4867 236
rect 4893 224 4899 256
rect 4877 124 4883 216
rect 4925 184 4931 256
rect 4941 184 4947 336
rect 4973 284 4979 536
rect 4989 324 4995 516
rect 5085 504 5091 597
rect 5133 584 5139 596
rect 5149 544 5155 616
rect 5229 584 5235 697
rect 5293 684 5299 956
rect 5309 884 5315 1216
rect 5389 1104 5395 1196
rect 5405 1144 5411 1156
rect 5469 924 5475 1316
rect 5533 1304 5539 1396
rect 5565 1384 5571 1456
rect 5581 1404 5587 1476
rect 5597 1384 5603 1476
rect 5549 1344 5555 1356
rect 5581 1324 5587 1376
rect 5629 1364 5635 1396
rect 5661 1364 5667 1476
rect 5693 1384 5699 1497
rect 5885 1484 5891 1496
rect 5773 1424 5779 1456
rect 5613 1244 5619 1356
rect 5725 1324 5731 1356
rect 5757 1324 5763 1376
rect 5789 1340 5795 1376
rect 5773 1324 5779 1336
rect 5693 1304 5699 1316
rect 5677 1264 5683 1276
rect 5709 1244 5715 1296
rect 5517 1164 5523 1236
rect 5533 1084 5539 1096
rect 5629 1064 5635 1136
rect 5485 924 5491 956
rect 5565 944 5571 1056
rect 5597 984 5603 1056
rect 5629 984 5635 1036
rect 5533 924 5539 936
rect 5421 704 5427 876
rect 5613 824 5619 936
rect 5645 904 5651 996
rect 5709 964 5715 1036
rect 5725 1004 5731 1116
rect 5757 1084 5763 1236
rect 5821 1204 5827 1476
rect 5837 1244 5843 1476
rect 5853 1384 5859 1436
rect 5901 1404 5907 1476
rect 5933 1384 5939 1476
rect 5949 1364 5955 1396
rect 5965 1384 5971 1396
rect 6045 1364 6051 1636
rect 6093 1504 6099 1836
rect 6125 1784 6131 1836
rect 6205 1724 6211 1876
rect 6253 1844 6259 2016
rect 6269 1944 6275 2036
rect 6285 1924 6291 1936
rect 6301 1884 6307 2036
rect 6413 1904 6419 1916
rect 6525 1904 6531 2096
rect 6589 2004 6595 2116
rect 6637 2044 6643 2136
rect 6653 2124 6659 2216
rect 6685 2184 6691 2296
rect 6701 2204 6707 2276
rect 6733 2244 6739 2276
rect 6749 2223 6755 2296
rect 6765 2284 6771 2356
rect 6861 2324 6867 2376
rect 6925 2364 6931 2676
rect 6941 2584 6947 2616
rect 6957 2584 6963 2636
rect 6973 2384 6979 2636
rect 6813 2244 6819 2316
rect 6861 2284 6867 2316
rect 6893 2284 6899 2296
rect 6909 2284 6915 2336
rect 6941 2304 6947 2316
rect 6733 2217 6755 2223
rect 6669 2064 6675 2136
rect 6685 2124 6691 2176
rect 6701 2144 6707 2176
rect 6733 2164 6739 2217
rect 6669 1984 6675 2036
rect 6317 1783 6323 1896
rect 6344 1806 6350 1814
rect 6358 1806 6364 1814
rect 6372 1806 6378 1814
rect 6386 1806 6392 1814
rect 6445 1784 6451 1856
rect 6461 1844 6467 1896
rect 6557 1884 6563 1936
rect 6596 1897 6611 1903
rect 6605 1864 6611 1897
rect 6717 1884 6723 2076
rect 6317 1777 6332 1783
rect 6445 1764 6451 1776
rect 6477 1764 6483 1836
rect 6109 1504 6115 1556
rect 6157 1524 6163 1596
rect 6173 1504 6179 1676
rect 5773 1064 5779 1116
rect 5789 1104 5795 1116
rect 5821 1084 5827 1196
rect 5869 1124 5875 1256
rect 5901 1124 5907 1156
rect 5949 1084 5955 1236
rect 5981 1104 5987 1136
rect 5853 1004 5859 1056
rect 5997 964 6003 1316
rect 6061 1224 6067 1436
rect 6109 1404 6115 1476
rect 6189 1464 6195 1476
rect 6205 1464 6211 1716
rect 6237 1584 6243 1716
rect 6333 1664 6339 1696
rect 6269 1504 6275 1616
rect 6221 1464 6227 1496
rect 6285 1484 6291 1516
rect 6381 1484 6387 1636
rect 6397 1564 6403 1756
rect 6445 1724 6451 1756
rect 6493 1744 6499 1856
rect 6525 1784 6531 1836
rect 6541 1744 6547 1756
rect 6573 1744 6579 1776
rect 6621 1764 6627 1856
rect 6589 1724 6595 1756
rect 6429 1584 6435 1656
rect 6461 1604 6467 1716
rect 6493 1704 6499 1716
rect 6589 1704 6595 1716
rect 6605 1704 6611 1736
rect 6621 1724 6627 1756
rect 6477 1604 6483 1696
rect 6637 1684 6643 1836
rect 6653 1664 6659 1856
rect 6701 1784 6707 1880
rect 6733 1864 6739 2156
rect 6749 2104 6755 2156
rect 6765 2124 6771 2236
rect 6781 2224 6787 2236
rect 6797 2144 6803 2156
rect 6829 2123 6835 2236
rect 6861 2144 6867 2276
rect 6909 2124 6915 2276
rect 6925 2164 6931 2216
rect 6989 2164 6995 2196
rect 6820 2117 6835 2123
rect 6749 1984 6755 2096
rect 6797 1984 6803 2116
rect 6781 1864 6787 1916
rect 6813 1864 6819 2056
rect 6877 1924 6883 1996
rect 6733 1844 6739 1856
rect 6797 1784 6803 1856
rect 6813 1804 6819 1856
rect 6845 1784 6851 1876
rect 6701 1763 6707 1776
rect 6685 1757 6707 1763
rect 6397 1524 6403 1556
rect 6125 1384 6131 1456
rect 6205 1403 6211 1436
rect 6189 1397 6211 1403
rect 6124 1350 6132 1356
rect 6189 1324 6195 1397
rect 6237 1344 6243 1456
rect 6344 1406 6350 1414
rect 6358 1406 6364 1414
rect 6372 1406 6378 1414
rect 6386 1406 6392 1414
rect 6029 1084 6035 1096
rect 6045 1043 6051 1076
rect 6020 1037 6051 1043
rect 5517 724 5523 816
rect 5693 704 5699 936
rect 5389 664 5395 676
rect 5437 664 5443 680
rect 5181 544 5187 556
rect 5156 537 5171 543
rect 5085 484 5091 496
rect 5101 384 5107 456
rect 5021 324 5027 356
rect 4989 304 4995 316
rect 4957 224 4963 256
rect 5021 144 5027 316
rect 5085 264 5091 276
rect 5101 144 5107 356
rect 5133 304 5139 336
rect 5165 324 5171 537
rect 5197 384 5203 536
rect 5261 504 5267 536
rect 5389 524 5395 656
rect 5453 564 5459 576
rect 5469 564 5475 636
rect 5485 544 5491 676
rect 5517 524 5523 636
rect 5565 604 5571 696
rect 5581 684 5587 696
rect 5197 324 5203 376
rect 5133 164 5139 176
rect 5149 164 5155 316
rect 5165 304 5171 316
rect 5197 264 5203 276
rect 5213 264 5219 496
rect 5229 344 5235 356
rect 5245 344 5251 476
rect 5181 124 5187 236
rect 5229 164 5235 216
rect 5053 104 5059 116
rect 5213 104 5219 136
rect 5245 104 5251 336
rect 5261 184 5267 496
rect 5309 284 5315 376
rect 5389 364 5395 516
rect 5565 504 5571 556
rect 5581 517 5596 523
rect 5421 384 5427 416
rect 5453 304 5459 396
rect 5340 264 5348 270
rect 5293 164 5299 196
rect 5341 144 5347 236
rect 5469 184 5475 276
rect 5485 264 5491 296
rect 5485 224 5491 256
rect 5533 144 5539 356
rect 5581 344 5587 517
rect 5597 504 5603 516
rect 5613 464 5619 536
rect 5629 343 5635 536
rect 5645 384 5651 694
rect 5709 584 5715 916
rect 5741 884 5747 956
rect 5997 943 6003 956
rect 6061 944 6067 1216
rect 6093 1064 6099 1096
rect 6109 1064 6115 1176
rect 6157 1104 6163 1296
rect 6173 1084 6179 1096
rect 6205 1084 6211 1196
rect 6221 1104 6227 1176
rect 6205 944 6211 1016
rect 6269 964 6275 976
rect 5981 937 6003 943
rect 5981 924 5987 937
rect 6285 924 6291 1376
rect 6413 1324 6419 1496
rect 6429 1244 6435 1576
rect 6541 1524 6547 1536
rect 6573 1504 6579 1636
rect 6445 1364 6451 1476
rect 6461 1384 6467 1456
rect 6557 1384 6563 1436
rect 6461 1344 6467 1356
rect 6573 1344 6579 1416
rect 6589 1364 6595 1656
rect 6621 1624 6627 1636
rect 6621 1464 6627 1496
rect 6653 1484 6659 1496
rect 6685 1444 6691 1757
rect 6733 1584 6739 1756
rect 6829 1744 6835 1756
rect 6749 1724 6755 1736
rect 6861 1704 6867 1876
rect 6877 1864 6883 1916
rect 6893 1904 6899 2036
rect 6925 2024 6931 2156
rect 7005 2144 7011 2356
rect 7037 2264 7043 2336
rect 7069 2284 7075 2676
rect 7117 2544 7123 2556
rect 7149 2544 7155 2716
rect 7181 2684 7187 2796
rect 7213 2704 7219 2716
rect 7325 2704 7331 2796
rect 7389 2784 7395 2936
rect 7357 2704 7363 2736
rect 7405 2704 7411 2716
rect 7453 2704 7459 2916
rect 7469 2904 7475 2916
rect 7485 2904 7491 2916
rect 7517 2884 7523 2956
rect 7661 2944 7667 2956
rect 7725 2944 7731 2996
rect 7773 2984 7779 3077
rect 7789 3044 7795 3076
rect 7485 2704 7491 2776
rect 7517 2704 7523 2716
rect 7549 2704 7555 2936
rect 7597 2924 7603 2936
rect 7629 2904 7635 2916
rect 7229 2544 7235 2636
rect 7245 2504 7251 2516
rect 7261 2503 7267 2696
rect 7373 2664 7379 2676
rect 7309 2644 7315 2656
rect 7277 2564 7283 2576
rect 7357 2544 7363 2556
rect 7252 2497 7267 2503
rect 7069 2144 7075 2156
rect 7101 2123 7107 2336
rect 7245 2324 7251 2496
rect 7117 2304 7123 2316
rect 7245 2304 7251 2316
rect 7229 2297 7244 2303
rect 7117 2144 7123 2176
rect 7133 2124 7139 2136
rect 7101 2117 7116 2123
rect 6957 2084 6963 2096
rect 7021 1924 7027 2036
rect 6893 1804 6899 1876
rect 6893 1764 6899 1776
rect 6925 1724 6931 1836
rect 6989 1784 6995 1856
rect 6781 1664 6787 1696
rect 6877 1684 6883 1716
rect 6877 1644 6883 1676
rect 7053 1584 7059 2116
rect 7069 2004 7075 2036
rect 7165 1983 7171 2276
rect 7181 2144 7187 2156
rect 7213 2144 7219 2176
rect 7229 2124 7235 2297
rect 7277 2284 7283 2456
rect 7357 2284 7363 2436
rect 7373 2304 7379 2656
rect 7389 2644 7395 2696
rect 7453 2664 7459 2676
rect 7469 2584 7475 2696
rect 7597 2684 7603 2696
rect 7661 2684 7667 2936
rect 7789 2924 7795 2956
rect 7837 2924 7843 2976
rect 7677 2684 7683 2696
rect 7485 2563 7491 2676
rect 7533 2664 7539 2676
rect 7469 2557 7491 2563
rect 7469 2384 7475 2557
rect 7485 2444 7491 2496
rect 7517 2484 7523 2596
rect 7565 2544 7571 2596
rect 7581 2584 7587 2656
rect 7645 2564 7651 2596
rect 7661 2564 7667 2676
rect 7677 2564 7683 2636
rect 7789 2624 7795 2916
rect 7805 2724 7811 2776
rect 7837 2704 7843 2856
rect 7837 2664 7843 2696
rect 7853 2684 7859 3276
rect 8013 3184 8019 3836
rect 8029 3263 8035 4196
rect 8045 4184 8051 4236
rect 8061 4144 8067 4396
rect 8077 4204 8083 4636
rect 8125 4624 8131 4676
rect 8141 4483 8147 5316
rect 8125 4477 8147 4483
rect 8093 4344 8099 4436
rect 8093 4144 8099 4296
rect 8045 3984 8051 4036
rect 8077 3924 8083 4136
rect 8093 4104 8099 4136
rect 8109 4124 8115 4236
rect 8093 4024 8099 4076
rect 8093 3984 8099 3996
rect 8109 3944 8115 3956
rect 8061 3864 8067 3916
rect 8109 3744 8115 3776
rect 8093 3584 8099 3716
rect 8045 3364 8051 3496
rect 8029 3257 8051 3263
rect 8029 3164 8035 3236
rect 7933 3124 7939 3136
rect 7869 3084 7875 3116
rect 8029 3104 8035 3116
rect 7908 3097 7923 3103
rect 7892 3077 7907 3083
rect 7869 2904 7875 3036
rect 7885 2784 7891 2876
rect 7901 2864 7907 3077
rect 7917 3064 7923 3097
rect 7933 2904 7939 2918
rect 7933 2784 7939 2856
rect 7869 2724 7875 2736
rect 7901 2684 7907 2736
rect 7949 2704 7955 3036
rect 7997 2724 8003 2916
rect 8013 2724 8019 2756
rect 7853 2644 7859 2676
rect 7917 2664 7923 2696
rect 7965 2664 7971 2696
rect 7549 2524 7555 2536
rect 7405 2304 7411 2316
rect 7149 1977 7171 1983
rect 7149 1884 7155 1977
rect 7197 1884 7203 1896
rect 7117 1764 7123 1836
rect 7213 1784 7219 2116
rect 7229 2104 7235 2116
rect 7261 2104 7267 2236
rect 7277 2204 7283 2276
rect 7293 2224 7299 2256
rect 7357 2224 7363 2256
rect 7293 2164 7299 2176
rect 7309 2124 7315 2196
rect 7373 2164 7379 2296
rect 7421 2264 7427 2376
rect 7501 2324 7507 2436
rect 7517 2384 7523 2476
rect 7469 2284 7475 2296
rect 7453 2264 7459 2276
rect 7517 2264 7523 2336
rect 7549 2304 7555 2516
rect 7581 2503 7587 2516
rect 7597 2503 7603 2556
rect 7581 2497 7603 2503
rect 7581 2324 7587 2497
rect 7613 2444 7619 2556
rect 7581 2264 7587 2316
rect 7597 2304 7603 2316
rect 7645 2284 7651 2556
rect 7684 2517 7699 2523
rect 7693 2324 7699 2517
rect 7741 2364 7747 2496
rect 7757 2343 7763 2496
rect 7789 2484 7795 2536
rect 7805 2524 7811 2536
rect 7821 2503 7827 2516
rect 7812 2497 7827 2503
rect 7748 2337 7763 2343
rect 7741 2304 7747 2336
rect 7773 2324 7779 2356
rect 7789 2324 7795 2476
rect 7757 2284 7763 2316
rect 7373 2144 7379 2156
rect 7325 1984 7331 2036
rect 7277 1904 7283 1976
rect 7357 1904 7363 2096
rect 7421 1923 7427 2136
rect 7421 1917 7443 1923
rect 7261 1784 7267 1796
rect 7181 1744 7187 1756
rect 7277 1744 7283 1896
rect 7325 1784 7331 1876
rect 7149 1644 7155 1736
rect 7341 1724 7347 1876
rect 7357 1724 7363 1896
rect 7437 1884 7443 1917
rect 7453 1904 7459 1916
rect 7469 1884 7475 2156
rect 7501 2144 7507 2236
rect 7789 2124 7795 2236
rect 7821 2144 7827 2296
rect 7837 2264 7843 2516
rect 7853 2304 7859 2636
rect 7805 2104 7811 2136
rect 7773 2084 7779 2096
rect 7805 1924 7811 1996
rect 7533 1884 7539 1896
rect 7597 1884 7603 1894
rect 7821 1884 7827 2136
rect 7869 2124 7875 2656
rect 7892 2537 7907 2543
rect 7901 2384 7907 2537
rect 8013 2524 8019 2636
rect 8029 2524 8035 3076
rect 8045 2684 8051 3257
rect 8061 3104 8067 3316
rect 8061 2984 8067 3076
rect 8077 2924 8083 3556
rect 8109 3324 8115 3716
rect 8109 3304 8115 3316
rect 8125 3283 8131 4477
rect 8141 4164 8147 4276
rect 8157 3724 8163 5636
rect 8109 3277 8131 3283
rect 8109 3023 8115 3277
rect 8093 3017 8115 3023
rect 8077 2584 8083 2916
rect 8093 2744 8099 3017
rect 8109 2604 8115 2636
rect 7917 2304 7923 2436
rect 8029 2304 8035 2516
rect 8109 2284 8115 2336
rect 7917 2264 7923 2276
rect 7949 2144 7955 2276
rect 7837 1884 7843 1916
rect 7853 1904 7859 2116
rect 7933 2084 7939 2118
rect 8061 2084 8067 2096
rect 8077 2083 8083 2116
rect 8068 2077 8083 2083
rect 7949 1924 7955 1936
rect 7965 1924 7971 1976
rect 8077 1904 8083 1936
rect 7812 1877 7820 1883
rect 7405 1784 7411 1856
rect 7373 1744 7379 1756
rect 7229 1684 7235 1716
rect 7357 1704 7363 1716
rect 7213 1664 7219 1676
rect 6749 1464 6755 1516
rect 6989 1504 6995 1536
rect 6893 1497 6908 1503
rect 6861 1484 6867 1496
rect 6877 1484 6883 1496
rect 6813 1464 6819 1476
rect 6749 1424 6755 1456
rect 6669 1384 6675 1396
rect 6589 1344 6595 1356
rect 6477 1284 6483 1316
rect 6317 1064 6323 1136
rect 6445 1104 6451 1236
rect 6509 1124 6515 1296
rect 6621 1264 6627 1296
rect 6637 1284 6643 1316
rect 6557 1184 6563 1236
rect 6477 1102 6483 1116
rect 6365 1084 6371 1096
rect 6301 1057 6316 1063
rect 6301 1024 6307 1057
rect 6317 963 6323 1036
rect 6344 1006 6350 1014
rect 6358 1006 6364 1014
rect 6372 1006 6378 1014
rect 6386 1006 6392 1014
rect 6445 964 6451 1076
rect 6461 964 6467 996
rect 6308 957 6323 963
rect 6301 924 6307 956
rect 5869 784 5875 896
rect 5741 544 5747 656
rect 5773 644 5779 656
rect 5805 644 5811 696
rect 5837 644 5843 656
rect 5853 623 5859 696
rect 5933 684 5939 816
rect 5949 724 5955 836
rect 5869 624 5875 676
rect 5901 664 5907 676
rect 5837 617 5859 623
rect 5805 584 5811 616
rect 5773 564 5779 576
rect 5837 564 5843 617
rect 5949 584 5955 716
rect 6141 702 6147 736
rect 6157 684 6163 916
rect 6237 904 6243 916
rect 6397 724 6403 956
rect 6477 944 6483 1036
rect 6573 944 6579 1096
rect 6589 1024 6595 1256
rect 6621 1144 6627 1236
rect 6653 1104 6659 1116
rect 6589 924 6595 1016
rect 6653 944 6659 1096
rect 6669 1084 6675 1236
rect 6685 1123 6691 1336
rect 6797 1324 6803 1336
rect 6701 1244 6707 1316
rect 6781 1204 6787 1316
rect 6749 1144 6755 1176
rect 6797 1143 6803 1316
rect 6813 1244 6819 1456
rect 6829 1284 6835 1476
rect 6893 1284 6899 1497
rect 6973 1344 6979 1476
rect 6781 1137 6803 1143
rect 6685 1117 6700 1123
rect 6733 1084 6739 1096
rect 6701 963 6707 1036
rect 6749 1023 6755 1116
rect 6765 1104 6771 1136
rect 6685 957 6707 963
rect 6733 1017 6755 1023
rect 6605 884 6611 936
rect 6685 924 6691 957
rect 6733 904 6739 1017
rect 6781 944 6787 1137
rect 6813 1044 6819 1116
rect 6829 1104 6835 1276
rect 6909 1263 6915 1336
rect 6925 1264 6931 1316
rect 6893 1257 6915 1263
rect 6893 1184 6899 1257
rect 6925 1144 6931 1236
rect 6973 1224 6979 1336
rect 6989 1304 6995 1476
rect 7005 1464 7011 1576
rect 7085 1524 7091 1556
rect 7181 1504 7187 1636
rect 7197 1604 7203 1636
rect 7261 1504 7267 1636
rect 7405 1584 7411 1636
rect 7437 1504 7443 1676
rect 7053 1404 7059 1496
rect 7117 1384 7123 1396
rect 7181 1324 7187 1496
rect 7085 1184 7091 1236
rect 7101 1184 7107 1296
rect 6845 1024 6851 1136
rect 7197 1124 7203 1416
rect 7309 1364 7315 1396
rect 7453 1344 7459 1736
rect 7613 1684 7619 1876
rect 7821 1726 7827 1836
rect 7917 1784 7923 1896
rect 7997 1864 8003 1876
rect 8045 1864 8051 1876
rect 7981 1764 7987 1836
rect 7501 1504 7507 1516
rect 7485 1484 7491 1496
rect 7549 1464 7555 1516
rect 7581 1504 7587 1656
rect 7645 1644 7651 1716
rect 7709 1584 7715 1718
rect 7805 1524 7811 1536
rect 7837 1497 7852 1503
rect 7533 1384 7539 1436
rect 7565 1343 7571 1436
rect 7597 1344 7603 1476
rect 7661 1464 7667 1476
rect 7645 1424 7651 1456
rect 7565 1337 7580 1343
rect 7677 1343 7683 1436
rect 7709 1424 7715 1496
rect 7677 1337 7692 1343
rect 7357 1324 7363 1336
rect 7405 1324 7411 1336
rect 7629 1324 7635 1336
rect 7693 1324 7699 1336
rect 7245 1284 7251 1318
rect 7533 1304 7539 1316
rect 7709 1304 7715 1356
rect 7245 1184 7251 1196
rect 7213 1124 7219 1136
rect 6957 1102 6963 1116
rect 7133 1084 7139 1096
rect 6877 1044 6883 1056
rect 6909 984 6915 1016
rect 7037 984 7043 1016
rect 7133 984 7139 1076
rect 7149 1044 7155 1076
rect 6893 964 6899 976
rect 7197 964 7203 1116
rect 7245 1104 7251 1116
rect 7277 1064 7283 1076
rect 7309 1024 7315 1116
rect 7325 1084 7331 1236
rect 7341 1184 7347 1276
rect 7645 1144 7651 1276
rect 7709 1164 7715 1296
rect 7373 1104 7379 1116
rect 7421 1084 7427 1096
rect 7437 1084 7443 1116
rect 7485 1084 7491 1096
rect 7421 1064 7427 1076
rect 7277 944 7283 996
rect 7357 944 7363 1036
rect 7373 944 7379 1036
rect 7012 937 7027 943
rect 6941 864 6947 936
rect 6973 904 6979 936
rect 7021 784 7027 937
rect 7053 904 7059 916
rect 7245 864 7251 918
rect 7117 764 7123 836
rect 6429 724 6435 736
rect 5821 544 5827 556
rect 5853 544 5859 556
rect 5613 337 5635 343
rect 5549 224 5555 256
rect 5581 184 5587 336
rect 5613 324 5619 337
rect 5597 304 5603 316
rect 5613 244 5619 316
rect 5629 304 5635 316
rect 5645 304 5651 336
rect 5677 324 5683 516
rect 5725 464 5731 536
rect 5741 524 5747 536
rect 5933 524 5939 556
rect 5693 384 5699 456
rect 5789 304 5795 516
rect 5837 324 5843 436
rect 5917 324 5923 456
rect 5629 264 5635 296
rect 5613 183 5619 236
rect 5597 177 5619 183
rect 5581 144 5587 176
rect 5597 144 5603 177
rect 5693 144 5699 296
rect 5725 284 5731 296
rect 5709 244 5715 256
rect 5789 244 5795 276
rect 5853 264 5859 316
rect 5901 284 5907 316
rect 5949 304 5955 576
rect 6013 544 6019 676
rect 6061 644 6067 656
rect 6077 543 6083 636
rect 6189 564 6195 696
rect 6333 684 6339 696
rect 6445 684 6451 696
rect 6477 684 6483 716
rect 6493 684 6499 736
rect 6317 644 6323 680
rect 6285 603 6291 636
rect 6344 606 6350 614
rect 6358 606 6364 614
rect 6372 606 6378 614
rect 6386 606 6392 614
rect 6269 597 6291 603
rect 6093 544 6099 556
rect 6068 537 6083 543
rect 5949 284 5955 296
rect 5853 164 5859 236
rect 5965 164 5971 516
rect 6157 484 6163 516
rect 6189 424 6195 556
rect 6237 544 6243 556
rect 6269 544 6275 597
rect 6285 524 6291 576
rect 6221 504 6227 516
rect 6253 324 6259 516
rect 6301 404 6307 556
rect 6333 524 6339 556
rect 6397 404 6403 516
rect 6413 504 6419 536
rect 6445 523 6451 556
rect 6461 544 6467 636
rect 6445 517 6460 523
rect 6477 484 6483 676
rect 6509 584 6515 636
rect 6509 524 6515 556
rect 6525 544 6531 696
rect 6541 583 6547 716
rect 6621 684 6627 696
rect 6541 577 6556 583
rect 6557 564 6563 576
rect 6525 504 6531 536
rect 6589 524 6595 656
rect 6605 544 6611 636
rect 6717 584 6723 676
rect 6749 664 6755 736
rect 6781 684 6787 696
rect 6813 624 6819 656
rect 6685 544 6691 576
rect 6765 544 6771 576
rect 6605 503 6611 536
rect 6669 504 6675 516
rect 6605 497 6620 503
rect 6484 477 6492 483
rect 6733 464 6739 516
rect 6749 504 6755 516
rect 6397 384 6403 396
rect 6445 384 6451 436
rect 6285 304 6291 376
rect 6701 304 6707 436
rect 6717 302 6723 356
rect 6237 284 6243 296
rect 6653 284 6659 296
rect 6813 284 6819 376
rect 6845 284 6851 676
rect 6861 584 6867 616
rect 6877 564 6883 596
rect 6941 564 6947 716
rect 7053 684 7059 696
rect 7213 684 7219 756
rect 7069 664 7075 676
rect 7277 664 7283 676
rect 7133 644 7139 656
rect 7021 544 7027 576
rect 7085 544 7091 636
rect 7133 563 7139 636
rect 7277 604 7283 656
rect 7197 564 7203 596
rect 7309 584 7315 896
rect 7341 884 7347 916
rect 7341 723 7347 836
rect 7373 724 7379 836
rect 7341 717 7356 723
rect 7325 684 7331 696
rect 7405 684 7411 896
rect 7421 764 7427 1056
rect 7437 1044 7443 1076
rect 7469 984 7475 1076
rect 7437 944 7443 976
rect 7485 924 7491 1076
rect 7549 1064 7555 1096
rect 7517 924 7523 936
rect 7549 904 7555 1016
rect 7565 984 7571 1076
rect 7597 944 7603 1136
rect 7613 1124 7619 1136
rect 7661 1104 7667 1116
rect 7677 1084 7683 1096
rect 7469 884 7475 896
rect 7469 784 7475 876
rect 7485 664 7491 716
rect 7517 684 7523 716
rect 7565 663 7571 916
rect 7629 884 7635 1036
rect 7677 684 7683 1076
rect 7725 1064 7731 1456
rect 7741 1304 7747 1476
rect 7757 1464 7763 1476
rect 7773 1444 7779 1496
rect 7757 1384 7763 1416
rect 7805 1344 7811 1456
rect 7821 1364 7827 1436
rect 7837 1384 7843 1497
rect 7869 1484 7875 1516
rect 7853 1344 7859 1476
rect 7901 1444 7907 1496
rect 7757 1304 7763 1316
rect 7837 1304 7843 1316
rect 7933 1304 7939 1436
rect 7981 1344 7987 1736
rect 8013 1726 8019 1756
rect 7997 1464 8003 1496
rect 8044 1464 8052 1470
rect 7757 1084 7763 1096
rect 7837 1084 7843 1296
rect 7885 1284 7891 1296
rect 7869 1104 7875 1236
rect 7933 1104 7939 1296
rect 7949 1284 7955 1316
rect 7981 1204 7987 1336
rect 7981 1104 7987 1136
rect 7853 1064 7859 1096
rect 7901 1084 7907 1096
rect 7556 657 7571 663
rect 7693 663 7699 1056
rect 7709 984 7715 1056
rect 7725 924 7731 1036
rect 7773 1024 7779 1056
rect 7789 1024 7795 1036
rect 7741 964 7747 996
rect 7805 944 7811 956
rect 7885 924 7891 1036
rect 7741 904 7747 918
rect 7997 904 8003 1036
rect 8013 964 8019 1196
rect 8029 1084 8035 1376
rect 8045 1344 8051 1436
rect 8061 1084 8067 1156
rect 8109 1084 8115 1496
rect 8061 1024 8067 1076
rect 8109 1064 8115 1076
rect 8013 944 8019 956
rect 8093 944 8099 1016
rect 8125 983 8131 2656
rect 8141 1924 8147 3096
rect 8157 2884 8163 2896
rect 8157 2084 8163 2096
rect 8141 1784 8147 1916
rect 8141 1164 8147 1236
rect 8157 1144 8163 1476
rect 8141 984 8147 1116
rect 8116 977 8131 983
rect 8109 940 8115 976
rect 8029 843 8035 918
rect 8029 837 8051 843
rect 7757 784 7763 836
rect 7773 664 7779 676
rect 7684 657 7699 663
rect 7117 557 7139 563
rect 7117 544 7123 557
rect 6973 517 6988 523
rect 6957 364 6963 436
rect 6973 384 6979 517
rect 6893 324 6899 336
rect 5933 144 5939 156
rect 5469 124 5475 136
rect 5709 124 5715 136
rect 5357 104 5363 116
rect 5725 104 5731 136
rect 5981 124 5987 236
rect 5885 104 5891 116
rect 6013 104 6019 276
rect 6093 124 6099 196
rect 6237 164 6243 276
rect 6317 257 6332 263
rect 6253 204 6259 236
rect 6109 144 6115 156
rect 6237 144 6243 156
rect 6285 124 6291 156
rect 5661 84 5667 96
rect 6317 84 6323 257
rect 6344 206 6350 214
rect 6358 206 6364 214
rect 6372 206 6378 214
rect 6386 206 6392 214
rect 6525 144 6531 156
rect 6589 144 6595 156
rect 6397 84 6403 116
rect 6461 104 6467 136
rect 6541 123 6547 136
rect 6573 124 6579 136
rect 6532 117 6547 123
rect 6605 104 6611 156
rect 6621 144 6627 256
rect 6781 204 6787 236
rect 6621 104 6627 136
rect 6653 104 6659 176
rect 6717 144 6723 196
rect 6813 184 6819 276
rect 6861 244 6867 276
rect 6733 164 6739 176
rect 6813 144 6819 156
rect 6829 124 6835 236
rect 6845 164 6851 236
rect 6877 144 6883 256
rect 6893 124 6899 276
rect 6925 264 6931 336
rect 6957 224 6963 336
rect 7037 323 7043 516
rect 7053 484 7059 516
rect 7085 504 7091 516
rect 7021 317 7043 323
rect 6973 284 6979 296
rect 6989 264 6995 316
rect 7005 244 7011 256
rect 6669 104 6675 116
rect 6925 104 6931 216
rect 6989 144 6995 196
rect 7005 124 7011 236
rect 7021 204 7027 317
rect 7069 304 7075 496
rect 7085 324 7091 356
rect 7117 344 7123 536
rect 7133 364 7139 536
rect 7357 524 7363 636
rect 7149 324 7155 436
rect 7053 284 7059 296
rect 7197 284 7203 336
rect 7037 264 7043 276
rect 7101 264 7107 276
rect 7213 224 7219 296
rect 7229 284 7235 296
rect 7245 263 7251 316
rect 7341 284 7347 516
rect 7245 257 7260 263
rect 7117 144 7123 176
rect 7341 164 7347 276
rect 7373 164 7379 596
rect 7469 584 7475 656
rect 7485 584 7491 656
rect 7469 383 7475 476
rect 7460 377 7475 383
rect 7501 324 7507 536
rect 7533 524 7539 636
rect 7677 564 7683 656
rect 7741 624 7747 656
rect 7581 524 7587 536
rect 7581 384 7587 516
rect 7693 304 7699 316
rect 7661 284 7667 296
rect 7629 244 7635 256
rect 7277 144 7283 156
rect 7581 144 7587 236
rect 7693 203 7699 236
rect 7693 197 7715 203
rect 7709 126 7715 197
rect 7757 184 7763 316
rect 7789 304 7795 396
rect 7805 304 7811 716
rect 7901 704 7907 836
rect 8045 784 8051 837
rect 8061 724 8067 736
rect 7981 684 7987 716
rect 8013 684 8019 696
rect 7837 644 7843 656
rect 7821 637 7836 643
rect 7805 284 7811 296
rect 7821 284 7827 637
rect 7853 324 7859 396
rect 7869 324 7875 676
rect 7917 624 7923 664
rect 7965 644 7971 676
rect 7933 544 7939 636
rect 7981 524 7987 636
rect 7997 504 8003 656
rect 8013 624 8019 676
rect 8029 664 8035 716
rect 8045 524 8051 696
rect 8061 564 8067 616
rect 8077 543 8083 736
rect 8093 684 8099 696
rect 8109 684 8115 696
rect 8093 584 8099 656
rect 8141 644 8147 836
rect 8157 664 8163 716
rect 8141 544 8147 636
rect 8068 537 8083 543
rect 8077 503 8083 537
rect 8125 504 8131 516
rect 8077 497 8092 503
rect 8061 484 8067 496
rect 7885 324 7891 436
rect 7917 404 7923 436
rect 7853 224 7859 236
rect 7869 204 7875 236
rect 7885 144 7891 316
rect 7917 304 7923 316
rect 8061 304 8067 476
rect 8093 304 8099 476
rect 7933 284 7939 296
rect 7229 104 7235 116
rect 7357 104 7363 116
rect 7917 104 7923 196
rect 7949 124 7955 236
rect 7965 224 7971 276
rect 8013 244 8019 296
rect 7965 144 7971 156
rect 7997 124 8003 176
rect 8013 144 8019 156
rect 8029 104 8035 276
rect 8045 144 8051 236
rect 8061 144 8067 296
rect 8077 164 8083 236
rect 8093 184 8099 236
rect 8093 124 8099 136
rect 7988 97 8012 103
rect 7357 84 7363 96
rect 8109 84 8115 396
rect 8157 284 8163 296
rect 1972 77 2003 83
rect 1736 6 1742 14
rect 1750 6 1756 14
rect 1764 6 1770 14
rect 1778 6 1784 14
rect 4808 6 4814 14
rect 4822 6 4828 14
rect 4836 6 4842 14
rect 4850 6 4856 14
<< m3contact >>
rect 684 5756 692 5764
rect 940 5756 948 5764
rect 988 5756 996 5764
rect 1036 5756 1044 5764
rect 1276 5756 1284 5764
rect 1484 5756 1492 5764
rect 2364 5756 2372 5764
rect 284 5736 292 5744
rect 332 5740 340 5744
rect 332 5736 340 5740
rect 92 5716 100 5724
rect 204 5716 212 5724
rect 236 5716 244 5724
rect 124 5696 132 5704
rect 76 5576 84 5584
rect 380 5716 388 5724
rect 364 5676 372 5684
rect 204 5656 212 5664
rect 364 5656 372 5664
rect 636 5736 644 5744
rect 508 5716 516 5724
rect 556 5696 564 5704
rect 860 5736 868 5744
rect 876 5736 884 5744
rect 700 5716 708 5724
rect 924 5716 932 5724
rect 748 5696 756 5704
rect 428 5676 436 5684
rect 540 5676 548 5684
rect 396 5556 404 5564
rect 252 5516 260 5524
rect 300 5516 308 5524
rect 204 5496 212 5504
rect 12 5376 20 5384
rect 332 5496 340 5504
rect 364 5496 372 5504
rect 220 5476 228 5484
rect 188 5456 196 5464
rect 268 5436 276 5444
rect 204 5376 212 5384
rect 140 5318 148 5324
rect 140 5316 148 5318
rect 220 5336 228 5344
rect 300 5476 308 5484
rect 348 5476 356 5484
rect 316 5456 324 5464
rect 300 5376 308 5384
rect 284 5336 292 5344
rect 316 5356 324 5364
rect 380 5476 388 5484
rect 492 5576 500 5584
rect 444 5556 452 5564
rect 428 5496 436 5504
rect 412 5476 420 5484
rect 476 5476 484 5484
rect 396 5456 404 5464
rect 428 5456 436 5464
rect 396 5436 404 5444
rect 412 5396 420 5404
rect 364 5356 372 5364
rect 316 5336 324 5344
rect 252 5316 260 5324
rect 268 5316 276 5324
rect 316 5316 324 5324
rect 396 5336 404 5344
rect 460 5436 468 5444
rect 460 5356 468 5364
rect 444 5316 452 5324
rect 348 5296 356 5304
rect 460 5296 468 5304
rect 428 5276 436 5284
rect 460 5276 468 5284
rect 716 5656 724 5664
rect 908 5676 916 5684
rect 508 5516 516 5524
rect 556 5516 564 5524
rect 908 5596 916 5604
rect 956 5596 964 5604
rect 1004 5716 1012 5724
rect 1036 5716 1044 5724
rect 1020 5656 1028 5664
rect 988 5556 996 5564
rect 972 5516 980 5524
rect 572 5496 580 5504
rect 972 5496 980 5504
rect 540 5396 548 5404
rect 604 5476 612 5484
rect 764 5476 772 5484
rect 620 5436 628 5444
rect 556 5376 564 5384
rect 572 5376 580 5384
rect 556 5356 564 5364
rect 636 5356 644 5364
rect 652 5356 660 5364
rect 620 5336 628 5344
rect 540 5316 548 5324
rect 524 5276 532 5284
rect 444 5256 452 5264
rect 204 5176 212 5184
rect 76 5096 84 5104
rect 204 5096 212 5104
rect 236 5096 244 5104
rect 268 5096 276 5104
rect 124 5056 132 5064
rect 204 5056 212 5064
rect 28 4956 36 4964
rect 188 5036 196 5044
rect 204 4996 212 5004
rect 140 4976 148 4984
rect 12 4936 20 4944
rect 44 4936 52 4944
rect 76 4916 84 4924
rect 188 4956 196 4964
rect 364 5076 372 5084
rect 556 5276 564 5284
rect 700 5356 708 5364
rect 716 5336 724 5344
rect 684 5316 692 5324
rect 1148 5736 1156 5744
rect 1484 5736 1492 5744
rect 1660 5736 1668 5744
rect 1868 5736 1876 5744
rect 2012 5736 2020 5744
rect 2204 5736 2212 5744
rect 1116 5716 1124 5724
rect 1164 5716 1172 5724
rect 1100 5676 1108 5684
rect 1196 5696 1204 5704
rect 1116 5656 1124 5664
rect 1068 5536 1076 5544
rect 1100 5536 1108 5544
rect 1148 5516 1156 5524
rect 1052 5496 1060 5504
rect 892 5456 900 5464
rect 940 5456 948 5464
rect 1052 5456 1060 5464
rect 876 5436 884 5444
rect 1036 5436 1044 5444
rect 844 5416 852 5424
rect 972 5416 980 5424
rect 1020 5416 1028 5424
rect 828 5376 836 5384
rect 844 5376 852 5384
rect 924 5376 932 5384
rect 940 5356 948 5364
rect 1132 5476 1140 5484
rect 1180 5676 1188 5684
rect 1180 5536 1188 5544
rect 1244 5676 1252 5684
rect 1244 5556 1252 5564
rect 1228 5516 1236 5524
rect 1228 5476 1236 5484
rect 1132 5456 1140 5464
rect 1164 5456 1172 5464
rect 1212 5416 1220 5424
rect 1324 5716 1332 5724
rect 1420 5718 1428 5724
rect 1420 5716 1428 5718
rect 1276 5696 1284 5704
rect 1324 5676 1332 5684
rect 1420 5696 1428 5704
rect 1580 5696 1588 5704
rect 1356 5676 1364 5684
rect 1340 5656 1348 5664
rect 1372 5536 1380 5544
rect 1340 5516 1348 5524
rect 1356 5496 1364 5504
rect 1212 5396 1220 5404
rect 1260 5396 1268 5404
rect 1100 5376 1108 5384
rect 1148 5376 1156 5384
rect 812 5316 820 5324
rect 844 5316 852 5324
rect 908 5316 916 5324
rect 668 5296 676 5304
rect 812 5296 820 5304
rect 668 5276 676 5284
rect 652 5256 660 5264
rect 604 5216 612 5224
rect 492 5096 500 5104
rect 604 5096 612 5104
rect 284 4996 292 5004
rect 252 4956 260 4964
rect 396 4976 404 4984
rect 316 4956 324 4964
rect 268 4936 276 4944
rect 268 4916 276 4924
rect 284 4916 292 4924
rect 172 4896 180 4904
rect 92 4876 100 4884
rect 156 4876 164 4884
rect 172 4776 180 4784
rect 140 4702 148 4704
rect 140 4696 148 4702
rect 220 4896 228 4904
rect 252 4896 260 4904
rect 188 4736 196 4744
rect 364 4936 372 4944
rect 428 4956 436 4964
rect 412 4936 420 4944
rect 348 4896 356 4904
rect 396 4896 404 4904
rect 380 4876 388 4884
rect 300 4836 308 4844
rect 284 4756 292 4764
rect 300 4736 308 4744
rect 268 4716 276 4724
rect 268 4696 276 4704
rect 220 4676 228 4684
rect 12 4636 20 4644
rect 204 4636 212 4644
rect 428 4876 436 4884
rect 412 4836 420 4844
rect 460 4996 468 5004
rect 460 4956 468 4964
rect 460 4916 468 4924
rect 460 4896 468 4904
rect 444 4816 452 4824
rect 364 4736 372 4744
rect 460 4736 468 4744
rect 348 4716 356 4724
rect 364 4696 372 4704
rect 396 4696 404 4704
rect 476 4716 484 4724
rect 252 4656 260 4664
rect 316 4656 324 4664
rect 252 4636 260 4644
rect 316 4576 324 4584
rect 348 4576 356 4584
rect 300 4556 308 4564
rect 236 4516 244 4524
rect 12 4396 20 4404
rect 28 4256 36 4264
rect 28 4236 36 4244
rect 108 4396 116 4404
rect 140 4356 148 4364
rect 172 4316 180 4324
rect 156 4276 164 4284
rect 108 4216 116 4224
rect 172 4156 180 4164
rect 412 4536 420 4544
rect 476 4536 484 4544
rect 364 4516 372 4524
rect 236 4336 244 4344
rect 220 4296 228 4304
rect 236 4276 244 4284
rect 300 4496 308 4504
rect 380 4496 388 4504
rect 412 4496 420 4504
rect 444 4516 452 4524
rect 300 4356 308 4364
rect 348 4356 356 4364
rect 284 4316 292 4324
rect 300 4316 308 4324
rect 348 4296 356 4304
rect 444 4476 452 4484
rect 428 4316 436 4324
rect 476 4296 484 4304
rect 380 4276 388 4284
rect 412 4276 420 4284
rect 236 4256 244 4264
rect 252 4256 260 4264
rect 204 4196 212 4204
rect 204 4156 212 4164
rect 140 4136 148 4144
rect 188 4136 196 4144
rect 252 4236 260 4244
rect 1292 5456 1300 5464
rect 1276 5376 1284 5384
rect 1308 5396 1316 5404
rect 1308 5376 1316 5384
rect 1244 5316 1252 5324
rect 1292 5316 1300 5324
rect 1132 5296 1140 5304
rect 1260 5296 1268 5304
rect 1292 5296 1300 5304
rect 1180 5196 1188 5204
rect 1116 5136 1124 5144
rect 1372 5316 1380 5324
rect 1468 5676 1476 5684
rect 1436 5496 1444 5504
rect 1452 5476 1460 5484
rect 1404 5436 1412 5444
rect 1548 5636 1556 5644
rect 1644 5696 1652 5704
rect 1612 5656 1620 5664
rect 1596 5576 1604 5584
rect 1628 5556 1636 5564
rect 1564 5536 1572 5544
rect 1612 5536 1620 5544
rect 1676 5696 1684 5704
rect 1548 5456 1556 5464
rect 1644 5456 1652 5464
rect 1660 5396 1668 5404
rect 1644 5376 1652 5384
rect 1500 5316 1508 5324
rect 1356 5296 1364 5304
rect 1356 5196 1364 5204
rect 1308 5156 1316 5164
rect 1276 5136 1284 5144
rect 1308 5136 1316 5144
rect 988 5096 996 5104
rect 1148 5096 1156 5104
rect 556 5056 564 5064
rect 524 5036 532 5044
rect 556 4956 564 4964
rect 556 4896 564 4904
rect 508 4876 516 4884
rect 524 4876 532 4884
rect 556 4856 564 4864
rect 524 4776 532 4784
rect 524 4556 532 4564
rect 508 4516 516 4524
rect 508 4476 516 4484
rect 588 5056 596 5064
rect 636 4976 644 4984
rect 780 4976 788 4984
rect 604 4916 612 4924
rect 636 4916 644 4924
rect 604 4896 612 4904
rect 636 4896 644 4904
rect 588 4876 596 4884
rect 652 4876 660 4884
rect 620 4816 628 4824
rect 588 4696 596 4704
rect 716 4896 724 4904
rect 748 4856 756 4864
rect 700 4836 708 4844
rect 684 4776 692 4784
rect 668 4736 676 4744
rect 652 4716 660 4724
rect 684 4716 692 4724
rect 716 4776 724 4784
rect 636 4696 644 4704
rect 764 4756 772 4764
rect 732 4696 740 4704
rect 652 4676 660 4684
rect 716 4676 724 4684
rect 604 4636 612 4644
rect 620 4636 628 4644
rect 588 4316 596 4324
rect 524 4296 532 4304
rect 572 4296 580 4304
rect 492 4256 500 4264
rect 508 4256 516 4264
rect 252 4216 260 4224
rect 332 4216 340 4224
rect 268 4196 276 4204
rect 364 4196 372 4204
rect 188 4116 196 4124
rect 60 4096 68 4104
rect 140 4096 148 4104
rect 76 4016 84 4024
rect 28 3896 36 3904
rect 92 3902 100 3904
rect 92 3896 100 3902
rect 204 3896 212 3904
rect 236 3896 244 3904
rect 28 3836 36 3844
rect 188 3776 196 3784
rect 428 4176 436 4184
rect 284 4116 292 4124
rect 540 4236 548 4244
rect 508 4216 516 4224
rect 492 4176 500 4184
rect 476 4136 484 4144
rect 828 4956 836 4964
rect 812 4936 820 4944
rect 812 4736 820 4744
rect 860 4936 868 4944
rect 1068 5076 1076 5084
rect 1132 5076 1140 5084
rect 1116 5056 1124 5064
rect 1100 5036 1108 5044
rect 1180 5036 1188 5044
rect 1148 4996 1156 5004
rect 1004 4956 1012 4964
rect 1244 5056 1252 5064
rect 1228 5036 1236 5044
rect 1260 4976 1268 4984
rect 1196 4956 1204 4964
rect 876 4916 884 4924
rect 1148 4916 1156 4924
rect 892 4876 900 4884
rect 844 4856 852 4864
rect 828 4716 836 4724
rect 876 4716 884 4724
rect 972 4716 980 4724
rect 1132 4716 1140 4724
rect 940 4676 948 4684
rect 860 4616 868 4624
rect 908 4616 916 4624
rect 1196 4916 1204 4924
rect 1260 4916 1268 4924
rect 1308 5096 1316 5104
rect 1308 5056 1316 5064
rect 1372 5096 1380 5104
rect 1612 5196 1620 5204
rect 1788 5716 1796 5724
rect 1820 5716 1828 5724
rect 1724 5696 1732 5704
rect 1788 5696 1796 5704
rect 1692 5676 1700 5684
rect 1788 5656 1796 5664
rect 1900 5676 1908 5684
rect 1836 5636 1844 5644
rect 1884 5636 1892 5644
rect 1742 5606 1750 5614
rect 1756 5606 1764 5614
rect 1770 5606 1778 5614
rect 1756 5456 1764 5464
rect 1852 5536 1860 5544
rect 1692 5356 1700 5364
rect 1740 5356 1748 5364
rect 1676 5336 1684 5344
rect 1708 5316 1716 5324
rect 1804 5416 1812 5424
rect 1756 5276 1764 5284
rect 1708 5216 1716 5224
rect 1742 5206 1750 5214
rect 1756 5206 1764 5214
rect 1770 5206 1778 5214
rect 1820 5396 1828 5404
rect 1868 5456 1876 5464
rect 2060 5716 2068 5724
rect 2252 5716 2260 5724
rect 2268 5716 2276 5724
rect 2380 5716 2388 5724
rect 1980 5656 1988 5664
rect 1980 5576 1988 5584
rect 1932 5556 1940 5564
rect 1996 5536 2004 5544
rect 2028 5536 2036 5544
rect 2092 5536 2100 5544
rect 2156 5536 2164 5544
rect 2220 5536 2228 5544
rect 1932 5496 1940 5504
rect 2028 5516 2036 5524
rect 1980 5496 1988 5504
rect 1948 5476 1956 5484
rect 1900 5436 1908 5444
rect 1964 5436 1972 5444
rect 2204 5516 2212 5524
rect 2092 5476 2100 5484
rect 2124 5476 2132 5484
rect 2172 5476 2180 5484
rect 1996 5456 2004 5464
rect 2028 5416 2036 5424
rect 2044 5396 2052 5404
rect 2044 5376 2052 5384
rect 2028 5356 2036 5364
rect 1916 5316 1924 5324
rect 1980 5316 1988 5324
rect 2028 5316 2036 5324
rect 1996 5276 2004 5284
rect 1916 5116 1924 5124
rect 2028 5096 2036 5104
rect 1340 5056 1348 5064
rect 1356 5036 1364 5044
rect 1308 4916 1316 4924
rect 1228 4896 1236 4904
rect 1404 5076 1412 5084
rect 1468 5076 1476 5084
rect 1516 5076 1524 5084
rect 1868 5076 1876 5084
rect 1548 4976 1556 4984
rect 1420 4956 1428 4964
rect 1324 4876 1332 4884
rect 1196 4776 1204 4784
rect 1356 4856 1364 4864
rect 1292 4776 1300 4784
rect 1308 4756 1316 4764
rect 1260 4716 1268 4724
rect 1180 4676 1188 4684
rect 1388 4716 1396 4724
rect 1292 4676 1300 4684
rect 1132 4656 1140 4664
rect 1260 4656 1268 4664
rect 1116 4636 1124 4644
rect 860 4596 868 4604
rect 972 4596 980 4604
rect 780 4576 788 4584
rect 812 4576 820 4584
rect 1004 4576 1012 4584
rect 1100 4576 1108 4584
rect 684 4518 692 4524
rect 684 4516 692 4518
rect 684 4496 692 4504
rect 700 4336 708 4344
rect 636 4316 644 4324
rect 684 4316 692 4324
rect 636 4276 644 4284
rect 636 4256 644 4264
rect 828 4516 836 4524
rect 892 4496 900 4504
rect 924 4396 932 4404
rect 780 4356 788 4364
rect 732 4316 740 4324
rect 732 4276 740 4284
rect 780 4276 788 4284
rect 828 4276 836 4284
rect 812 4256 820 4264
rect 876 4176 884 4184
rect 908 4156 916 4164
rect 988 4516 996 4524
rect 956 4396 964 4404
rect 988 4356 996 4364
rect 972 4296 980 4304
rect 1068 4516 1076 4524
rect 1132 4518 1140 4524
rect 1132 4516 1140 4518
rect 1020 4496 1028 4504
rect 1164 4496 1172 4504
rect 1052 4476 1060 4484
rect 1084 4476 1092 4484
rect 1036 4456 1044 4464
rect 1132 4456 1140 4464
rect 1148 4356 1156 4364
rect 1020 4316 1028 4324
rect 1052 4316 1060 4324
rect 1100 4296 1108 4304
rect 1052 4276 1060 4284
rect 1036 4256 1044 4264
rect 1004 4176 1012 4184
rect 1052 4156 1060 4164
rect 716 4136 724 4144
rect 892 4136 900 4144
rect 940 4136 948 4144
rect 956 4136 964 4144
rect 684 4116 692 4124
rect 748 4118 756 4124
rect 748 4116 756 4118
rect 588 4096 596 4104
rect 636 4096 644 4104
rect 540 4056 548 4064
rect 316 4016 324 4024
rect 444 4016 452 4024
rect 476 4016 484 4024
rect 540 3956 548 3964
rect 284 3936 292 3944
rect 412 3902 420 3904
rect 412 3896 420 3902
rect 220 3836 228 3844
rect 204 3756 212 3764
rect 124 3736 132 3744
rect 12 3516 20 3524
rect 76 3516 84 3524
rect 60 3476 68 3484
rect 44 3456 52 3464
rect 140 3476 148 3484
rect 188 3516 196 3524
rect 316 3736 324 3744
rect 284 3716 292 3724
rect 492 3836 500 3844
rect 492 3716 500 3724
rect 268 3696 276 3704
rect 348 3696 356 3704
rect 460 3696 468 3704
rect 412 3596 420 3604
rect 268 3516 276 3524
rect 492 3676 500 3684
rect 476 3636 484 3644
rect 220 3496 228 3504
rect 332 3496 340 3504
rect 460 3496 468 3504
rect 492 3516 500 3524
rect 380 3476 388 3484
rect 140 3456 148 3464
rect 236 3456 244 3464
rect 316 3456 324 3464
rect 364 3456 372 3464
rect 108 3436 116 3444
rect 76 3336 84 3344
rect 44 3276 52 3284
rect 140 3296 148 3304
rect 92 3116 100 3124
rect 12 3056 20 3064
rect 236 3436 244 3444
rect 236 3356 244 3364
rect 172 3336 180 3344
rect 76 3096 84 3104
rect 140 3096 148 3104
rect 188 3316 196 3324
rect 252 3336 260 3344
rect 348 3316 356 3324
rect 204 3296 212 3304
rect 284 3276 292 3284
rect 476 3456 484 3464
rect 572 3936 580 3944
rect 556 3896 564 3904
rect 524 3856 532 3864
rect 684 4036 692 4044
rect 732 4036 740 4044
rect 636 3916 644 3924
rect 588 3816 596 3824
rect 668 3896 676 3904
rect 780 3916 788 3924
rect 844 3916 852 3924
rect 780 3896 788 3904
rect 812 3896 820 3904
rect 844 3896 852 3904
rect 716 3876 724 3884
rect 684 3856 692 3864
rect 668 3816 676 3824
rect 540 3736 548 3744
rect 572 3736 580 3744
rect 652 3736 660 3744
rect 700 3776 708 3784
rect 764 3776 772 3784
rect 716 3736 724 3744
rect 828 3816 836 3824
rect 700 3716 708 3724
rect 716 3716 724 3724
rect 764 3656 772 3664
rect 1004 4096 1012 4104
rect 1260 4356 1268 4364
rect 1228 4296 1236 4304
rect 1132 4276 1140 4284
rect 1180 4276 1188 4284
rect 1196 4276 1204 4284
rect 1244 4276 1252 4284
rect 1116 4256 1124 4264
rect 1132 4196 1140 4204
rect 1100 4136 1108 4144
rect 1036 4116 1044 4124
rect 1068 4096 1076 4104
rect 1244 4156 1252 4164
rect 1116 4116 1124 4124
rect 1164 4116 1172 4124
rect 1116 4096 1124 4104
rect 1148 4096 1156 4104
rect 1084 4076 1092 4084
rect 1164 4076 1172 4084
rect 1148 4056 1156 4064
rect 924 4036 932 4044
rect 1020 4036 1028 4044
rect 1084 4036 1092 4044
rect 940 3956 948 3964
rect 876 3896 884 3904
rect 892 3876 900 3884
rect 1004 3876 1012 3884
rect 1052 3876 1060 3884
rect 860 3856 868 3864
rect 1020 3856 1028 3864
rect 908 3816 916 3824
rect 1036 3816 1044 3824
rect 860 3796 868 3804
rect 892 3796 900 3804
rect 972 3776 980 3784
rect 860 3736 868 3744
rect 924 3736 932 3744
rect 956 3736 964 3744
rect 1020 3756 1028 3764
rect 988 3736 996 3744
rect 1036 3736 1044 3744
rect 1068 3776 1076 3784
rect 1068 3756 1076 3764
rect 1100 3936 1108 3944
rect 1260 4036 1268 4044
rect 1212 3916 1220 3924
rect 1292 4296 1300 4304
rect 1292 4256 1300 4264
rect 1100 3876 1108 3884
rect 1148 3876 1156 3884
rect 1116 3736 1124 3744
rect 892 3716 900 3724
rect 1052 3716 1060 3724
rect 1116 3696 1124 3704
rect 908 3676 916 3684
rect 972 3676 980 3684
rect 1100 3676 1108 3684
rect 812 3656 820 3664
rect 796 3616 804 3624
rect 572 3596 580 3604
rect 396 3376 404 3384
rect 396 3356 404 3364
rect 444 3336 452 3344
rect 460 3336 468 3344
rect 396 3316 404 3324
rect 428 3316 436 3324
rect 428 3296 436 3304
rect 460 3296 468 3304
rect 236 3116 244 3124
rect 380 3116 388 3124
rect 60 3076 68 3084
rect 108 3076 116 3084
rect 156 3076 164 3084
rect 60 3056 68 3064
rect 92 3036 100 3044
rect 28 2936 36 2944
rect 60 2936 68 2944
rect 44 2916 52 2924
rect 28 2896 36 2904
rect 44 2856 52 2864
rect 76 2856 84 2864
rect 172 3056 180 3064
rect 284 3076 292 3084
rect 188 3036 196 3044
rect 140 2936 148 2944
rect 188 2936 196 2944
rect 220 2936 228 2944
rect 300 2936 308 2944
rect 204 2916 212 2924
rect 140 2896 148 2904
rect 172 2896 180 2904
rect 204 2896 212 2904
rect 508 3436 516 3444
rect 940 3616 948 3624
rect 668 3496 676 3504
rect 860 3496 868 3504
rect 540 3476 548 3484
rect 492 3416 500 3424
rect 524 3416 532 3424
rect 508 3396 516 3404
rect 572 3336 580 3344
rect 540 3316 548 3324
rect 604 3316 612 3324
rect 492 3296 500 3304
rect 588 3296 596 3304
rect 524 3276 532 3284
rect 524 3156 532 3164
rect 476 3136 484 3144
rect 492 3116 500 3124
rect 540 3136 548 3144
rect 412 3076 420 3084
rect 524 3076 532 3084
rect 604 3216 612 3224
rect 636 3476 644 3484
rect 1004 3536 1012 3544
rect 1020 3496 1028 3504
rect 1004 3476 1012 3484
rect 924 3436 932 3444
rect 956 3436 964 3444
rect 732 3396 740 3404
rect 796 3396 804 3404
rect 636 3336 644 3344
rect 700 3336 708 3344
rect 684 3316 692 3324
rect 668 3256 676 3264
rect 620 3196 628 3204
rect 636 3176 644 3184
rect 668 3156 676 3164
rect 700 3256 708 3264
rect 572 3116 580 3124
rect 732 3316 740 3324
rect 764 3316 772 3324
rect 892 3336 900 3344
rect 828 3316 836 3324
rect 892 3316 900 3324
rect 988 3316 996 3324
rect 780 3276 788 3284
rect 748 3256 756 3264
rect 716 3236 724 3244
rect 748 3236 756 3244
rect 732 3196 740 3204
rect 700 3136 708 3144
rect 652 3076 660 3084
rect 732 3076 740 3084
rect 428 3036 436 3044
rect 460 2996 468 3004
rect 364 2956 372 2964
rect 188 2856 196 2864
rect 364 2856 372 2864
rect 204 2776 212 2784
rect 236 2776 244 2784
rect 268 2736 276 2744
rect 396 2736 404 2744
rect 156 2716 164 2724
rect 316 2716 324 2724
rect 428 2716 436 2724
rect 124 2696 132 2704
rect 268 2696 276 2704
rect 108 2676 116 2684
rect 556 3056 564 3064
rect 636 3056 644 3064
rect 716 3056 724 3064
rect 556 2996 564 3004
rect 556 2976 564 2984
rect 620 2976 628 2984
rect 492 2936 500 2944
rect 588 2936 596 2944
rect 684 3036 692 3044
rect 764 3216 772 3224
rect 780 3136 788 3144
rect 764 3116 772 3124
rect 956 3276 964 3284
rect 940 3256 948 3264
rect 1132 3576 1140 3584
rect 1100 3556 1108 3564
rect 1052 3496 1060 3504
rect 1116 3456 1124 3464
rect 1196 3856 1204 3864
rect 1244 3836 1252 3844
rect 1260 3836 1268 3844
rect 1324 4656 1332 4664
rect 1388 4656 1396 4664
rect 1452 4916 1460 4924
rect 1580 4956 1588 4964
rect 1500 4916 1508 4924
rect 1436 4896 1444 4904
rect 1580 4916 1588 4924
rect 1612 4936 1620 4944
rect 1516 4896 1524 4904
rect 1468 4856 1476 4864
rect 1452 4796 1460 4804
rect 1484 4796 1492 4804
rect 1436 4736 1444 4744
rect 1484 4716 1492 4724
rect 1452 4676 1460 4684
rect 1500 4676 1508 4684
rect 1532 4656 1540 4664
rect 1324 4596 1332 4604
rect 1420 4596 1428 4604
rect 1548 4596 1556 4604
rect 1532 4556 1540 4564
rect 1340 4436 1348 4444
rect 1356 4356 1364 4364
rect 1324 4256 1332 4264
rect 1388 4436 1396 4444
rect 1596 4876 1604 4884
rect 2092 5336 2100 5344
rect 2140 5456 2148 5464
rect 2172 5336 2180 5344
rect 2220 5496 2228 5504
rect 2252 5496 2260 5504
rect 2204 5356 2212 5364
rect 2332 5696 2340 5704
rect 2380 5696 2388 5704
rect 2412 5676 2420 5684
rect 2348 5516 2356 5524
rect 2300 5456 2308 5464
rect 2300 5436 2308 5444
rect 2236 5336 2244 5344
rect 2284 5336 2292 5344
rect 2252 5316 2260 5324
rect 2076 5296 2084 5304
rect 2108 5276 2116 5284
rect 2460 5756 2468 5764
rect 2588 5756 2596 5764
rect 2492 5696 2500 5704
rect 2476 5676 2484 5684
rect 3278 5806 3286 5814
rect 3292 5806 3300 5814
rect 3306 5806 3314 5814
rect 2812 5796 2820 5804
rect 2844 5796 2852 5804
rect 3020 5796 3028 5804
rect 3068 5796 3076 5804
rect 3612 5796 3620 5804
rect 3644 5796 3652 5804
rect 2732 5776 2740 5784
rect 2828 5776 2836 5784
rect 2604 5736 2612 5744
rect 2652 5736 2660 5744
rect 2572 5716 2580 5724
rect 2620 5696 2628 5704
rect 2636 5676 2644 5684
rect 2444 5656 2452 5664
rect 2540 5656 2548 5664
rect 2700 5716 2708 5724
rect 2812 5716 2820 5724
rect 2668 5656 2676 5664
rect 2812 5696 2820 5704
rect 2716 5676 2724 5684
rect 2780 5676 2788 5684
rect 2700 5576 2708 5584
rect 2668 5536 2676 5544
rect 2540 5516 2548 5524
rect 2828 5656 2836 5664
rect 2796 5576 2804 5584
rect 2428 5496 2436 5504
rect 2476 5496 2484 5504
rect 2668 5496 2676 5504
rect 2444 5476 2452 5484
rect 2492 5476 2500 5484
rect 2380 5396 2388 5404
rect 2412 5356 2420 5364
rect 2620 5356 2628 5364
rect 2444 5336 2452 5344
rect 2604 5336 2612 5344
rect 2332 5316 2340 5324
rect 2268 5276 2276 5284
rect 2220 5256 2228 5264
rect 2380 5316 2388 5324
rect 2476 5318 2484 5324
rect 2476 5316 2484 5318
rect 2396 5296 2404 5304
rect 2668 5336 2676 5344
rect 2988 5736 2996 5744
rect 3148 5776 3156 5784
rect 3292 5776 3300 5784
rect 2924 5716 2932 5724
rect 3036 5696 3044 5704
rect 3052 5676 3060 5684
rect 3084 5656 3092 5664
rect 3084 5596 3092 5604
rect 3356 5736 3364 5744
rect 3548 5736 3556 5744
rect 3276 5716 3284 5724
rect 3404 5716 3412 5724
rect 3452 5716 3460 5724
rect 3596 5716 3604 5724
rect 3228 5696 3236 5704
rect 3196 5676 3204 5684
rect 3148 5596 3156 5604
rect 3116 5576 3124 5584
rect 2908 5536 2916 5544
rect 2860 5516 2868 5524
rect 3532 5696 3540 5704
rect 3532 5676 3540 5684
rect 3628 5676 3636 5684
rect 3628 5656 3636 5664
rect 3596 5576 3604 5584
rect 3436 5516 3444 5524
rect 3548 5516 3556 5524
rect 2844 5496 2852 5504
rect 2940 5496 2948 5504
rect 3004 5502 3012 5504
rect 3004 5496 3012 5502
rect 3324 5496 3332 5504
rect 3436 5496 3444 5504
rect 3468 5496 3476 5504
rect 3532 5496 3540 5504
rect 3564 5496 3572 5504
rect 3676 5756 3684 5764
rect 3884 5756 3892 5764
rect 3948 5756 3956 5764
rect 3740 5736 3748 5744
rect 3868 5736 3876 5744
rect 3676 5716 3684 5724
rect 3644 5496 3652 5504
rect 3724 5696 3732 5704
rect 3772 5696 3780 5704
rect 6350 5806 6358 5814
rect 6364 5806 6372 5814
rect 6378 5806 6386 5814
rect 6156 5796 6164 5804
rect 6204 5796 6212 5804
rect 4508 5776 4516 5784
rect 4764 5776 4772 5784
rect 5020 5776 5028 5784
rect 6140 5776 6148 5784
rect 4156 5756 4164 5764
rect 3964 5736 3972 5744
rect 3836 5676 3844 5684
rect 3772 5496 3780 5504
rect 2892 5476 2900 5484
rect 3036 5476 3044 5484
rect 3420 5476 3428 5484
rect 3516 5476 3524 5484
rect 3580 5476 3588 5484
rect 2940 5456 2948 5464
rect 2764 5396 2772 5404
rect 2828 5396 2836 5404
rect 2844 5376 2852 5384
rect 3100 5456 3108 5464
rect 3132 5416 3140 5424
rect 3900 5596 3908 5604
rect 4092 5716 4100 5724
rect 4284 5716 4292 5724
rect 4060 5696 4068 5704
rect 4108 5696 4116 5704
rect 3996 5676 4004 5684
rect 3996 5636 4004 5644
rect 4044 5636 4052 5644
rect 4012 5616 4020 5624
rect 3964 5576 3972 5584
rect 3916 5496 3924 5504
rect 3980 5502 3988 5504
rect 3980 5496 3988 5502
rect 4332 5636 4340 5644
rect 4204 5616 4212 5624
rect 4092 5596 4100 5604
rect 4108 5596 4116 5604
rect 4172 5596 4180 5604
rect 4268 5596 4276 5604
rect 4044 5496 4052 5504
rect 4108 5576 4116 5584
rect 4124 5516 4132 5524
rect 3916 5476 3924 5484
rect 4076 5476 4084 5484
rect 4092 5476 4100 5484
rect 3628 5456 3636 5464
rect 3708 5456 3716 5464
rect 3836 5456 3844 5464
rect 3228 5416 3236 5424
rect 3278 5406 3286 5414
rect 3292 5406 3300 5414
rect 3306 5406 3314 5414
rect 3500 5376 3508 5384
rect 3100 5356 3108 5364
rect 3132 5356 3140 5364
rect 3164 5356 3172 5364
rect 3356 5356 3364 5364
rect 2908 5336 2916 5344
rect 3004 5336 3012 5344
rect 3052 5336 3060 5344
rect 3084 5336 3092 5344
rect 2860 5316 2868 5324
rect 2892 5318 2900 5324
rect 2892 5316 2900 5318
rect 3068 5316 3076 5324
rect 3164 5336 3172 5344
rect 3052 5296 3060 5304
rect 2604 5276 2612 5284
rect 2636 5276 2644 5284
rect 2364 5256 2372 5264
rect 2140 5176 2148 5184
rect 2348 5176 2356 5184
rect 2220 5136 2228 5144
rect 2332 5136 2340 5144
rect 2540 5136 2548 5144
rect 2748 5136 2756 5144
rect 2188 5116 2196 5124
rect 2236 5116 2244 5124
rect 2444 5116 2452 5124
rect 2460 5116 2468 5124
rect 2492 5116 2500 5124
rect 2556 5116 2564 5124
rect 2620 5116 2628 5124
rect 2668 5116 2676 5124
rect 2732 5116 2740 5124
rect 2428 5096 2436 5104
rect 2156 5076 2164 5084
rect 2236 5076 2244 5084
rect 2252 5076 2260 5084
rect 2268 5076 2276 5084
rect 2140 5056 2148 5064
rect 1804 4936 1812 4944
rect 1932 4936 1940 4944
rect 1964 4936 1972 4944
rect 2012 4876 2020 4884
rect 1724 4836 1732 4844
rect 1980 4836 1988 4844
rect 1742 4806 1750 4814
rect 1756 4806 1764 4814
rect 1770 4806 1778 4814
rect 1644 4776 1652 4784
rect 1628 4756 1636 4764
rect 1820 4736 1828 4744
rect 1820 4716 1828 4724
rect 1580 4676 1588 4684
rect 1628 4676 1636 4684
rect 1852 4696 1860 4704
rect 2124 4956 2132 4964
rect 2092 4896 2100 4904
rect 2140 4896 2148 4904
rect 2140 4876 2148 4884
rect 2188 5056 2196 5064
rect 2220 4956 2228 4964
rect 2300 4996 2308 5004
rect 2348 4936 2356 4944
rect 2364 4936 2372 4944
rect 2396 4936 2404 4944
rect 2428 4936 2436 4944
rect 2444 4936 2452 4944
rect 2236 4916 2244 4924
rect 2300 4916 2308 4924
rect 2172 4896 2180 4904
rect 2220 4896 2228 4904
rect 2444 4916 2452 4924
rect 2572 5096 2580 5104
rect 2476 5076 2484 5084
rect 2524 5076 2532 5084
rect 2588 5076 2596 5084
rect 2604 5076 2612 5084
rect 2668 5076 2676 5084
rect 2492 4956 2500 4964
rect 2668 5056 2676 5064
rect 2700 5056 2708 5064
rect 2572 4996 2580 5004
rect 2588 4976 2596 4984
rect 2540 4936 2548 4944
rect 2668 4956 2676 4964
rect 2636 4936 2644 4944
rect 2684 4936 2692 4944
rect 2732 4936 2740 4944
rect 3020 5216 3028 5224
rect 2860 5136 2868 5144
rect 2924 5116 2932 5124
rect 2956 5116 2964 5124
rect 2876 5076 2884 5084
rect 3180 5316 3188 5324
rect 3516 5356 3524 5364
rect 3532 5336 3540 5344
rect 3580 5336 3588 5344
rect 3324 5296 3332 5304
rect 3564 5316 3572 5324
rect 3708 5416 3716 5424
rect 3836 5416 3844 5424
rect 3644 5336 3652 5344
rect 3692 5336 3700 5344
rect 3212 5256 3220 5264
rect 3484 5256 3492 5264
rect 3548 5256 3556 5264
rect 3116 5216 3124 5224
rect 3164 5216 3172 5224
rect 3100 5096 3108 5104
rect 3004 5076 3012 5084
rect 2956 5056 2964 5064
rect 3004 5016 3012 5024
rect 2924 4996 2932 5004
rect 2908 4976 2916 4984
rect 3052 5016 3060 5024
rect 3100 4976 3108 4984
rect 3212 5136 3220 5144
rect 3244 5116 3252 5124
rect 3356 5116 3364 5124
rect 3212 5076 3220 5084
rect 3212 4996 3220 5004
rect 2796 4936 2804 4944
rect 2812 4936 2820 4944
rect 2892 4936 2900 4944
rect 3020 4936 3028 4944
rect 3228 4976 3236 4984
rect 3340 5096 3348 5104
rect 3468 5096 3476 5104
rect 3372 5076 3380 5084
rect 3340 5056 3348 5064
rect 3278 5006 3286 5014
rect 3292 5006 3300 5014
rect 3306 5006 3314 5014
rect 3228 4956 3236 4964
rect 3324 4956 3332 4964
rect 3340 4956 3348 4964
rect 2524 4916 2532 4924
rect 2572 4916 2580 4924
rect 2636 4916 2644 4924
rect 2700 4916 2708 4924
rect 2300 4896 2308 4904
rect 2332 4896 2340 4904
rect 2380 4896 2388 4904
rect 2652 4896 2660 4904
rect 2764 4896 2772 4904
rect 2780 4896 2788 4904
rect 2828 4896 2836 4904
rect 2860 4896 2868 4904
rect 3148 4916 3156 4924
rect 2972 4896 2980 4904
rect 3180 4896 3188 4904
rect 2172 4876 2180 4884
rect 2252 4876 2260 4884
rect 2396 4876 2404 4884
rect 2460 4876 2468 4884
rect 2524 4876 2532 4884
rect 2876 4876 2884 4884
rect 3212 4876 3220 4884
rect 2156 4856 2164 4864
rect 2380 4856 2388 4864
rect 3148 4856 3156 4864
rect 3196 4836 3204 4844
rect 2092 4796 2100 4804
rect 2572 4796 2580 4804
rect 2668 4796 2676 4804
rect 2236 4776 2244 4784
rect 2044 4756 2052 4764
rect 2044 4736 2052 4744
rect 2124 4736 2132 4744
rect 2108 4716 2116 4724
rect 1708 4656 1716 4664
rect 1596 4556 1604 4564
rect 1612 4556 1620 4564
rect 1580 4536 1588 4544
rect 1580 4516 1588 4524
rect 1900 4676 1908 4684
rect 1804 4576 1812 4584
rect 1852 4576 1860 4584
rect 1740 4556 1748 4564
rect 1692 4536 1700 4544
rect 1676 4516 1684 4524
rect 1740 4516 1748 4524
rect 1820 4516 1828 4524
rect 1500 4496 1508 4504
rect 1612 4496 1620 4504
rect 1742 4406 1750 4414
rect 1756 4406 1764 4414
rect 1770 4406 1778 4414
rect 1404 4316 1412 4324
rect 1500 4316 1508 4324
rect 1660 4316 1668 4324
rect 1436 4296 1444 4304
rect 1548 4296 1556 4304
rect 1708 4296 1716 4304
rect 1772 4302 1780 4304
rect 1772 4296 1780 4302
rect 1404 4256 1412 4264
rect 1388 4196 1396 4204
rect 1356 4116 1364 4124
rect 1372 4116 1380 4124
rect 1324 3976 1332 3984
rect 1388 3916 1396 3924
rect 1452 4276 1460 4284
rect 1532 4276 1540 4284
rect 1532 4256 1540 4264
rect 1436 4176 1444 4184
rect 1452 4156 1460 4164
rect 1516 4156 1524 4164
rect 1436 4136 1444 4144
rect 1500 4136 1508 4144
rect 1612 4276 1620 4284
rect 1628 4256 1636 4264
rect 1708 4256 1716 4264
rect 1580 4156 1588 4164
rect 1596 4136 1604 4144
rect 1500 4116 1508 4124
rect 1724 4156 1732 4164
rect 1756 4156 1764 4164
rect 1612 4116 1620 4124
rect 1628 4116 1636 4124
rect 1564 4096 1572 4104
rect 1644 4096 1652 4104
rect 1420 4076 1428 4084
rect 1532 4056 1540 4064
rect 1420 3976 1428 3984
rect 1742 4006 1750 4014
rect 1756 4006 1764 4014
rect 1770 4006 1778 4014
rect 1692 3936 1700 3944
rect 1580 3916 1588 3924
rect 1628 3916 1636 3924
rect 1516 3896 1524 3904
rect 1308 3876 1316 3884
rect 1452 3876 1460 3884
rect 1292 3796 1300 3804
rect 1356 3856 1364 3864
rect 1340 3816 1348 3824
rect 1468 3816 1476 3824
rect 1276 3756 1284 3764
rect 1212 3696 1220 3704
rect 1244 3676 1252 3684
rect 1228 3516 1236 3524
rect 1180 3496 1188 3504
rect 1228 3496 1236 3504
rect 1164 3456 1172 3464
rect 1228 3396 1236 3404
rect 1148 3376 1156 3384
rect 1228 3376 1236 3384
rect 1292 3556 1300 3564
rect 1436 3796 1444 3804
rect 1516 3796 1524 3804
rect 1836 4296 1844 4304
rect 1868 4256 1876 4264
rect 1868 4236 1876 4244
rect 1836 4176 1844 4184
rect 1852 4176 1860 4184
rect 1820 4136 1828 4144
rect 1916 4596 1924 4604
rect 2124 4696 2132 4704
rect 2076 4676 2084 4684
rect 2108 4676 2116 4684
rect 2060 4596 2068 4604
rect 2092 4636 2100 4644
rect 2172 4696 2180 4704
rect 2460 4756 2468 4764
rect 2284 4736 2292 4744
rect 2412 4716 2420 4724
rect 2364 4696 2372 4704
rect 2444 4696 2452 4704
rect 2220 4676 2228 4684
rect 2156 4656 2164 4664
rect 2140 4636 2148 4644
rect 1980 4516 1988 4524
rect 2204 4516 2212 4524
rect 2124 4496 2132 4504
rect 2252 4656 2260 4664
rect 2300 4636 2308 4644
rect 2380 4636 2388 4644
rect 2428 4656 2436 4664
rect 2412 4556 2420 4564
rect 2364 4536 2372 4544
rect 2396 4536 2404 4544
rect 2268 4518 2276 4524
rect 2268 4516 2276 4518
rect 2220 4476 2228 4484
rect 1996 4456 2004 4464
rect 2044 4456 2052 4464
rect 2108 4436 2116 4444
rect 1916 4316 1924 4324
rect 2076 4336 2084 4344
rect 2092 4316 2100 4324
rect 1964 4236 1972 4244
rect 1996 4276 2004 4284
rect 1980 4216 1988 4224
rect 1900 4176 1908 4184
rect 1916 4156 1924 4164
rect 2012 4156 2020 4164
rect 1932 4136 1940 4144
rect 1900 4096 1908 4104
rect 1932 4096 1940 4104
rect 2076 4276 2084 4284
rect 2204 4336 2212 4344
rect 2236 4336 2244 4344
rect 2268 4336 2276 4344
rect 2156 4316 2164 4324
rect 2140 4256 2148 4264
rect 2108 4196 2116 4204
rect 2156 4236 2164 4244
rect 2028 4136 2036 4144
rect 2140 4136 2148 4144
rect 2044 4116 2052 4124
rect 2252 4256 2260 4264
rect 2204 4236 2212 4244
rect 2476 4696 2484 4704
rect 2524 4696 2532 4704
rect 2460 4676 2468 4684
rect 2492 4656 2500 4664
rect 2476 4596 2484 4604
rect 2332 4516 2340 4524
rect 2444 4516 2452 4524
rect 2364 4496 2372 4504
rect 2460 4496 2468 4504
rect 2348 4476 2356 4484
rect 2540 4556 2548 4564
rect 2492 4516 2500 4524
rect 2524 4516 2532 4524
rect 2540 4496 2548 4504
rect 2412 4476 2420 4484
rect 2444 4476 2452 4484
rect 2540 4476 2548 4484
rect 2380 4456 2388 4464
rect 2396 4316 2404 4324
rect 2316 4296 2324 4304
rect 2460 4296 2468 4304
rect 2556 4296 2564 4304
rect 2268 4156 2276 4164
rect 2316 4136 2324 4144
rect 2188 4116 2196 4124
rect 2236 4116 2244 4124
rect 2188 4096 2196 4104
rect 1996 4056 2004 4064
rect 1884 4036 1892 4044
rect 1868 3916 1876 3924
rect 1932 3936 1940 3944
rect 1628 3896 1636 3904
rect 1756 3896 1764 3904
rect 1804 3896 1812 3904
rect 1900 3896 1908 3904
rect 1964 3896 1972 3904
rect 2092 3896 2100 3904
rect 1660 3856 1668 3864
rect 1484 3736 1492 3744
rect 1532 3736 1540 3744
rect 1708 3756 1716 3764
rect 1852 3856 1860 3864
rect 1836 3836 1844 3844
rect 1964 3876 1972 3884
rect 2044 3876 2052 3884
rect 1884 3856 1892 3864
rect 1916 3856 1924 3864
rect 1820 3816 1828 3824
rect 1740 3756 1748 3764
rect 1644 3736 1652 3744
rect 1724 3736 1732 3744
rect 1804 3736 1812 3744
rect 1532 3716 1540 3724
rect 1612 3716 1620 3724
rect 1372 3556 1380 3564
rect 1356 3536 1364 3544
rect 1404 3536 1412 3544
rect 1260 3516 1268 3524
rect 1308 3496 1316 3504
rect 1452 3576 1460 3584
rect 1436 3516 1444 3524
rect 1372 3496 1380 3504
rect 1436 3496 1444 3504
rect 1580 3696 1588 3704
rect 1676 3696 1684 3704
rect 1516 3656 1524 3664
rect 1548 3656 1556 3664
rect 1660 3656 1668 3664
rect 1724 3656 1732 3664
rect 1516 3556 1524 3564
rect 1484 3536 1492 3544
rect 1500 3536 1508 3544
rect 1612 3536 1620 3544
rect 1628 3516 1636 3524
rect 1564 3496 1572 3504
rect 1340 3476 1348 3484
rect 1548 3476 1556 3484
rect 1820 3716 1828 3724
rect 1820 3676 1828 3684
rect 1804 3636 1812 3644
rect 1742 3606 1750 3614
rect 1756 3606 1764 3614
rect 1770 3606 1778 3614
rect 1644 3496 1652 3504
rect 1676 3496 1684 3504
rect 1676 3476 1684 3484
rect 1420 3456 1428 3464
rect 1596 3456 1604 3464
rect 1708 3456 1716 3464
rect 1324 3416 1332 3424
rect 1324 3376 1332 3384
rect 1036 3356 1044 3364
rect 1068 3316 1076 3324
rect 1020 3296 1028 3304
rect 1004 3236 1012 3244
rect 924 3216 932 3224
rect 844 3196 852 3204
rect 1132 3318 1140 3324
rect 1132 3316 1140 3318
rect 1100 3296 1108 3304
rect 1036 3276 1044 3284
rect 1068 3196 1076 3204
rect 1052 3156 1060 3164
rect 828 3116 836 3124
rect 1004 3096 1012 3104
rect 828 3076 836 3084
rect 892 3076 900 3084
rect 908 3076 916 3084
rect 956 3076 964 3084
rect 764 3056 772 3064
rect 796 2976 804 2984
rect 780 2936 788 2944
rect 748 2876 756 2884
rect 748 2856 756 2864
rect 732 2836 740 2844
rect 508 2756 516 2764
rect 844 3036 852 3044
rect 828 2956 836 2964
rect 812 2876 820 2884
rect 780 2836 788 2844
rect 1740 3416 1748 3424
rect 1612 3396 1620 3404
rect 1788 3396 1796 3404
rect 1484 3356 1492 3364
rect 1308 3316 1316 3324
rect 1276 3156 1284 3164
rect 1276 3136 1284 3144
rect 1148 3096 1156 3104
rect 1180 3096 1188 3104
rect 1148 3076 1156 3084
rect 1212 3076 1220 3084
rect 1276 3076 1284 3084
rect 1164 3036 1172 3044
rect 1004 2996 1012 3004
rect 924 2940 932 2944
rect 924 2936 932 2940
rect 876 2876 884 2884
rect 604 2716 612 2724
rect 620 2716 628 2724
rect 492 2696 500 2704
rect 572 2696 580 2704
rect 428 2676 436 2684
rect 476 2636 484 2644
rect 476 2596 484 2604
rect 140 2536 148 2544
rect 604 2676 612 2684
rect 540 2576 548 2584
rect 588 2576 596 2584
rect 508 2556 516 2564
rect 540 2556 548 2564
rect 508 2496 516 2504
rect 108 2276 116 2284
rect 76 2196 84 2204
rect 300 2356 308 2364
rect 204 2316 212 2324
rect 188 2236 196 2244
rect 220 2236 228 2244
rect 156 2216 164 2224
rect 188 2216 196 2224
rect 156 2196 164 2204
rect 188 2156 196 2164
rect 124 2136 132 2144
rect 268 2236 276 2244
rect 236 2196 244 2204
rect 204 2136 212 2144
rect 220 2136 228 2144
rect 476 2396 484 2404
rect 364 2356 372 2364
rect 300 2236 308 2244
rect 108 2116 116 2124
rect 140 2116 148 2124
rect 172 2116 180 2124
rect 204 2096 212 2104
rect 12 2076 20 2084
rect 76 2076 84 2084
rect 28 1896 36 1904
rect 60 1902 68 1904
rect 60 1896 68 1902
rect 252 2116 260 2124
rect 284 2196 292 2204
rect 252 2076 260 2084
rect 220 1956 228 1964
rect 204 1916 212 1924
rect 348 2336 356 2344
rect 380 2316 388 2324
rect 444 2316 452 2324
rect 348 2276 356 2284
rect 508 2356 516 2364
rect 508 2316 516 2324
rect 540 2316 548 2324
rect 412 2276 420 2284
rect 476 2276 484 2284
rect 364 2196 372 2204
rect 396 2196 404 2204
rect 572 2396 580 2404
rect 492 2156 500 2164
rect 828 2696 836 2704
rect 892 2696 900 2704
rect 956 2736 964 2744
rect 876 2676 884 2684
rect 940 2676 948 2684
rect 988 2676 996 2684
rect 764 2656 772 2664
rect 732 2636 740 2644
rect 620 2536 628 2544
rect 796 2656 804 2664
rect 844 2656 852 2664
rect 924 2636 932 2644
rect 940 2576 948 2584
rect 796 2556 804 2564
rect 908 2556 916 2564
rect 924 2556 932 2564
rect 732 2456 740 2464
rect 604 2356 612 2364
rect 652 2316 660 2324
rect 604 2296 612 2304
rect 620 2196 628 2204
rect 524 2136 532 2144
rect 300 2116 308 2124
rect 460 2116 468 2124
rect 572 2116 580 2124
rect 348 2096 356 2104
rect 636 2136 644 2144
rect 892 2536 900 2544
rect 812 2516 820 2524
rect 844 2516 852 2524
rect 860 2516 868 2524
rect 892 2516 900 2524
rect 940 2496 948 2504
rect 892 2476 900 2484
rect 844 2436 852 2444
rect 780 2376 788 2384
rect 844 2376 852 2384
rect 764 2296 772 2304
rect 1132 2956 1140 2964
rect 1084 2936 1092 2944
rect 1164 2936 1172 2944
rect 1260 2976 1268 2984
rect 1244 2856 1252 2864
rect 1052 2716 1060 2724
rect 1068 2696 1076 2704
rect 1164 2716 1172 2724
rect 1116 2696 1124 2704
rect 1100 2676 1108 2684
rect 1020 2656 1028 2664
rect 1036 2596 1044 2604
rect 988 2556 996 2564
rect 1004 2536 1012 2544
rect 1084 2536 1092 2544
rect 972 2516 980 2524
rect 1036 2516 1044 2524
rect 1020 2496 1028 2504
rect 1100 2496 1108 2504
rect 1068 2476 1076 2484
rect 1532 3336 1540 3344
rect 1724 3336 1732 3344
rect 1756 3336 1764 3344
rect 1484 3296 1492 3304
rect 1356 3216 1364 3224
rect 1580 3276 1588 3284
rect 1532 3236 1540 3244
rect 1660 3296 1668 3304
rect 1612 3276 1620 3284
rect 1628 3276 1636 3284
rect 1676 3276 1684 3284
rect 1612 3236 1620 3244
rect 1596 3216 1604 3224
rect 1742 3206 1750 3214
rect 1756 3206 1764 3214
rect 1770 3206 1778 3214
rect 1900 3736 1908 3744
rect 2012 3856 2020 3864
rect 2092 3856 2100 3864
rect 2012 3756 2020 3764
rect 1868 3716 1876 3724
rect 1932 3716 1940 3724
rect 1964 3718 1972 3724
rect 1964 3716 1972 3718
rect 1836 3616 1844 3624
rect 2028 3736 2036 3744
rect 2140 3756 2148 3764
rect 2108 3736 2116 3744
rect 2156 3736 2164 3744
rect 2092 3716 2100 3724
rect 2140 3716 2148 3724
rect 2220 3756 2228 3764
rect 2316 4056 2324 4064
rect 2268 3996 2276 4004
rect 2396 4256 2404 4264
rect 2588 4736 2596 4744
rect 2588 4716 2596 4724
rect 3132 4776 3140 4784
rect 2860 4756 2868 4764
rect 2732 4736 2740 4744
rect 2828 4736 2836 4744
rect 2796 4716 2804 4724
rect 2844 4716 2852 4724
rect 3052 4716 3060 4724
rect 3116 4716 3124 4724
rect 2764 4696 2772 4704
rect 2796 4676 2804 4684
rect 2588 4636 2596 4644
rect 2812 4596 2820 4604
rect 2684 4556 2692 4564
rect 2764 4556 2772 4564
rect 2716 4536 2724 4544
rect 2748 4516 2756 4524
rect 2924 4696 2932 4704
rect 2972 4676 2980 4684
rect 3068 4656 3076 4664
rect 2828 4556 2836 4564
rect 2860 4556 2868 4564
rect 3164 4796 3172 4804
rect 3196 4716 3204 4724
rect 3180 4676 3188 4684
rect 3164 4656 3172 4664
rect 3228 4676 3236 4684
rect 3420 5076 3428 5084
rect 3452 5076 3460 5084
rect 3548 5216 3556 5224
rect 3676 5316 3684 5324
rect 4220 5496 4228 5504
rect 4332 5516 4340 5524
rect 4284 5476 4292 5484
rect 4252 5456 4260 5464
rect 4012 5396 4020 5404
rect 4060 5396 4068 5404
rect 3772 5356 3780 5364
rect 3868 5356 3876 5364
rect 3916 5356 3924 5364
rect 4028 5356 4036 5364
rect 3884 5316 3892 5324
rect 3660 5256 3668 5264
rect 3596 5196 3604 5204
rect 3516 5136 3524 5144
rect 3516 5116 3524 5124
rect 3548 5116 3556 5124
rect 3628 5116 3636 5124
rect 3484 5056 3492 5064
rect 3500 5056 3508 5064
rect 3388 4976 3396 4984
rect 3388 4956 3396 4964
rect 3420 4956 3428 4964
rect 3356 4916 3364 4924
rect 3372 4916 3380 4924
rect 3500 4936 3508 4944
rect 3420 4876 3428 4884
rect 3644 5096 3652 5104
rect 3548 5076 3556 5084
rect 3580 5076 3588 5084
rect 3580 5056 3588 5064
rect 3612 5056 3620 5064
rect 3660 5056 3668 5064
rect 3564 4996 3572 5004
rect 3644 4996 3652 5004
rect 3580 4936 3588 4944
rect 3612 4936 3620 4944
rect 3564 4916 3572 4924
rect 3548 4896 3556 4904
rect 3484 4876 3492 4884
rect 3532 4876 3540 4884
rect 3404 4856 3412 4864
rect 3468 4856 3476 4864
rect 3356 4696 3364 4704
rect 3548 4776 3556 4784
rect 3596 4736 3604 4744
rect 3628 4736 3636 4744
rect 3596 4716 3604 4724
rect 3420 4702 3428 4704
rect 3420 4696 3428 4702
rect 3516 4696 3524 4704
rect 3404 4676 3412 4684
rect 3276 4636 3284 4644
rect 3244 4616 3252 4624
rect 3278 4606 3286 4614
rect 3292 4606 3300 4614
rect 3306 4606 3314 4614
rect 3228 4576 3236 4584
rect 3244 4576 3252 4584
rect 3292 4576 3300 4584
rect 3324 4556 3332 4564
rect 2876 4536 2884 4544
rect 2972 4536 2980 4544
rect 3084 4536 3092 4544
rect 3148 4536 3156 4544
rect 3180 4536 3188 4544
rect 3212 4536 3220 4544
rect 3244 4536 3252 4544
rect 2860 4516 2868 4524
rect 2652 4496 2660 4504
rect 2684 4496 2692 4504
rect 2716 4496 2724 4504
rect 2796 4496 2804 4504
rect 2908 4496 2916 4504
rect 2924 4496 2932 4504
rect 3036 4496 3044 4504
rect 2668 4476 2676 4484
rect 2796 4476 2804 4484
rect 2812 4356 2820 4364
rect 3004 4356 3012 4364
rect 2700 4336 2708 4344
rect 2492 4276 2500 4284
rect 2412 4216 2420 4224
rect 2460 4256 2468 4264
rect 2428 4196 2436 4204
rect 2588 4216 2596 4224
rect 2540 4196 2548 4204
rect 2908 4336 2916 4344
rect 2876 4316 2884 4324
rect 2940 4316 2948 4324
rect 3228 4476 3236 4484
rect 3196 4436 3204 4444
rect 3260 4436 3268 4444
rect 2780 4296 2788 4304
rect 2844 4296 2852 4304
rect 2988 4296 2996 4304
rect 3020 4296 3028 4304
rect 2684 4256 2692 4264
rect 2716 4276 2724 4284
rect 2764 4276 2772 4284
rect 2812 4276 2820 4284
rect 2716 4236 2724 4244
rect 2700 4196 2708 4204
rect 2620 4156 2628 4164
rect 2684 4156 2692 4164
rect 2476 4136 2484 4144
rect 2444 4116 2452 4124
rect 2508 4116 2516 4124
rect 2364 4096 2372 4104
rect 2332 4016 2340 4024
rect 2380 4016 2388 4024
rect 2412 3936 2420 3944
rect 2444 3976 2452 3984
rect 2428 3916 2436 3924
rect 2284 3896 2292 3904
rect 2348 3896 2356 3904
rect 2300 3876 2308 3884
rect 2252 3816 2260 3824
rect 2460 3876 2468 3884
rect 2444 3856 2452 3864
rect 2268 3756 2276 3764
rect 2236 3736 2244 3744
rect 2284 3736 2292 3744
rect 2460 3776 2468 3784
rect 2316 3756 2324 3764
rect 2396 3756 2404 3764
rect 2380 3716 2388 3724
rect 2588 4116 2596 4124
rect 2524 4016 2532 4024
rect 2540 3956 2548 3964
rect 2524 3936 2532 3944
rect 2508 3916 2516 3924
rect 2572 3956 2580 3964
rect 2556 3916 2564 3924
rect 2604 4016 2612 4024
rect 2572 3856 2580 3864
rect 2508 3756 2516 3764
rect 2604 3856 2612 3864
rect 2604 3736 2612 3744
rect 2460 3716 2468 3724
rect 2476 3716 2484 3724
rect 2556 3716 2564 3724
rect 2220 3696 2228 3704
rect 2252 3696 2260 3704
rect 2348 3696 2356 3704
rect 2396 3696 2404 3704
rect 2444 3696 2452 3704
rect 2316 3576 2324 3584
rect 2396 3576 2404 3584
rect 2316 3556 2324 3564
rect 1852 3536 1860 3544
rect 1836 3376 1844 3384
rect 1804 3196 1812 3204
rect 1356 3136 1364 3144
rect 1404 3136 1412 3144
rect 1436 3136 1444 3144
rect 1340 3116 1348 3124
rect 1372 3116 1380 3124
rect 1340 3096 1348 3104
rect 1420 3096 1428 3104
rect 1372 3076 1380 3084
rect 1564 3116 1572 3124
rect 1644 3116 1652 3124
rect 1532 3096 1540 3104
rect 1580 3096 1588 3104
rect 1516 3076 1524 3084
rect 1388 3056 1396 3064
rect 1500 3056 1508 3064
rect 1612 3056 1620 3064
rect 1356 3036 1364 3044
rect 1324 2996 1332 3004
rect 1324 2976 1332 2984
rect 1404 2996 1412 3004
rect 1564 2996 1572 3004
rect 1660 3096 1668 3104
rect 1884 3516 1892 3524
rect 2156 3516 2164 3524
rect 2268 3516 2276 3524
rect 2268 3496 2276 3504
rect 2348 3516 2356 3524
rect 2636 4116 2644 4124
rect 2668 4116 2676 4124
rect 2716 4116 2724 4124
rect 2700 4096 2708 4104
rect 2636 3996 2644 4004
rect 2700 3956 2708 3964
rect 2684 3936 2692 3944
rect 2668 3916 2676 3924
rect 2828 4236 2836 4244
rect 3068 4276 3076 4284
rect 3020 4256 3028 4264
rect 3052 4256 3060 4264
rect 3020 4236 3028 4244
rect 2924 4216 2932 4224
rect 2876 4196 2884 4204
rect 2924 4196 2932 4204
rect 2908 4156 2916 4164
rect 2780 4116 2788 4124
rect 2812 4116 2820 4124
rect 2764 4096 2772 4104
rect 2780 4096 2788 4104
rect 2796 4096 2804 4104
rect 2780 4016 2788 4024
rect 2764 3996 2772 4004
rect 2732 3936 2740 3944
rect 2700 3916 2708 3924
rect 2732 3916 2740 3924
rect 2636 3876 2644 3884
rect 2684 3876 2692 3884
rect 2732 3876 2740 3884
rect 2780 3876 2788 3884
rect 2700 3856 2708 3864
rect 2732 3856 2740 3864
rect 2748 3796 2756 3804
rect 2796 3856 2804 3864
rect 2796 3836 2804 3844
rect 2652 3736 2660 3744
rect 2684 3736 2692 3744
rect 2684 3716 2692 3724
rect 2780 3696 2788 3704
rect 2908 4096 2916 4104
rect 2876 4076 2884 4084
rect 2828 3876 2836 3884
rect 2828 3856 2836 3864
rect 2844 3796 2852 3804
rect 2860 3796 2868 3804
rect 2844 3756 2852 3764
rect 2812 3716 2820 3724
rect 3148 4236 3156 4244
rect 3052 4216 3060 4224
rect 3116 4216 3124 4224
rect 2988 4156 2996 4164
rect 2956 4116 2964 4124
rect 2972 4096 2980 4104
rect 2940 4076 2948 4084
rect 2988 3996 2996 4004
rect 3084 4096 3092 4104
rect 3132 3976 3140 3984
rect 3260 4256 3268 4264
rect 3564 4696 3572 4704
rect 3564 4676 3572 4684
rect 3532 4656 3540 4664
rect 3580 4656 3588 4664
rect 3692 4996 3700 5004
rect 3676 4916 3684 4924
rect 3804 5156 3812 5164
rect 3756 5136 3764 5144
rect 3788 5136 3796 5144
rect 3724 5116 3732 5124
rect 3788 5116 3796 5124
rect 3724 5096 3732 5104
rect 3740 5076 3748 5084
rect 3852 5116 3860 5124
rect 4092 5336 4100 5344
rect 4172 5416 4180 5424
rect 4204 5376 4212 5384
rect 4156 5336 4164 5344
rect 4220 5336 4228 5344
rect 3948 5316 3956 5324
rect 4012 5316 4020 5324
rect 4140 5316 4148 5324
rect 4188 5316 4196 5324
rect 4268 5396 4276 5404
rect 4332 5456 4340 5464
rect 4332 5416 4340 5424
rect 4300 5376 4308 5384
rect 4396 5736 4404 5744
rect 4460 5716 4468 5724
rect 4556 5756 4564 5764
rect 4588 5756 4596 5764
rect 4524 5716 4532 5724
rect 4556 5716 4564 5724
rect 4492 5676 4500 5684
rect 4508 5676 4516 5684
rect 4380 5596 4388 5604
rect 4380 5556 4388 5564
rect 4620 5718 4628 5724
rect 4620 5716 4628 5718
rect 4684 5716 4692 5724
rect 4620 5636 4628 5644
rect 4988 5736 4996 5744
rect 4844 5716 4852 5724
rect 4732 5576 4740 5584
rect 4412 5556 4420 5564
rect 4588 5556 4596 5564
rect 4396 5536 4404 5544
rect 4380 5516 4388 5524
rect 4364 5496 4372 5504
rect 4572 5536 4580 5544
rect 4524 5516 4532 5524
rect 4556 5516 4564 5524
rect 4444 5496 4452 5504
rect 4460 5456 4468 5464
rect 4284 5336 4292 5344
rect 4348 5336 4356 5344
rect 4236 5316 4244 5324
rect 4252 5316 4260 5324
rect 3980 5296 3988 5304
rect 4220 5296 4228 5304
rect 4268 5296 4276 5304
rect 3900 5196 3908 5204
rect 3900 5096 3908 5104
rect 3884 5076 3892 5084
rect 3836 5056 3844 5064
rect 3740 4976 3748 4984
rect 3820 4976 3828 4984
rect 3708 4876 3716 4884
rect 3676 4856 3684 4864
rect 3804 4876 3812 4884
rect 3820 4876 3828 4884
rect 3708 4776 3716 4784
rect 3692 4716 3700 4724
rect 3724 4736 3732 4744
rect 3772 4736 3780 4744
rect 3980 5256 3988 5264
rect 3932 5076 3940 5084
rect 3884 5036 3892 5044
rect 3916 5036 3924 5044
rect 3900 5016 3908 5024
rect 3868 4916 3876 4924
rect 3836 4796 3844 4804
rect 3820 4756 3828 4764
rect 3644 4676 3652 4684
rect 3772 4676 3780 4684
rect 3676 4656 3684 4664
rect 3756 4656 3764 4664
rect 3692 4616 3700 4624
rect 3724 4596 3732 4604
rect 3564 4556 3572 4564
rect 3644 4556 3652 4564
rect 3404 4496 3412 4504
rect 3436 4476 3444 4484
rect 3516 4476 3524 4484
rect 3420 4316 3428 4324
rect 3452 4296 3460 4304
rect 3532 4296 3540 4304
rect 3324 4256 3332 4264
rect 3292 4236 3300 4244
rect 3278 4206 3286 4214
rect 3292 4206 3300 4214
rect 3306 4206 3314 4214
rect 3212 4196 3220 4204
rect 3180 4176 3188 4184
rect 3436 4276 3444 4284
rect 3436 4256 3444 4264
rect 3388 4176 3396 4184
rect 3356 4156 3364 4164
rect 3180 4136 3188 4144
rect 3340 4136 3348 4144
rect 3372 4136 3380 4144
rect 3468 4136 3476 4144
rect 3324 4116 3332 4124
rect 3196 4096 3204 4104
rect 3164 3936 3172 3944
rect 2956 3916 2964 3924
rect 3148 3916 3156 3924
rect 3212 3956 3220 3964
rect 3324 4016 3332 4024
rect 3308 3916 3316 3924
rect 3180 3896 3188 3904
rect 2956 3876 2964 3884
rect 2972 3876 2980 3884
rect 3052 3876 3060 3884
rect 2924 3856 2932 3864
rect 2908 3836 2916 3844
rect 2924 3836 2932 3844
rect 2940 3796 2948 3804
rect 3004 3856 3012 3864
rect 3052 3856 3060 3864
rect 3116 3856 3124 3864
rect 3148 3856 3156 3864
rect 3036 3796 3044 3804
rect 3148 3816 3156 3824
rect 3532 4276 3540 4284
rect 3580 4516 3588 4524
rect 3612 4516 3620 4524
rect 3884 4896 3892 4904
rect 3868 4696 3876 4704
rect 4012 5136 4020 5144
rect 3980 5096 3988 5104
rect 4540 5476 4548 5484
rect 4620 5476 4628 5484
rect 4556 5456 4564 5464
rect 4492 5416 4500 5424
rect 4748 5416 4756 5424
rect 4814 5606 4822 5614
rect 4828 5606 4836 5614
rect 4842 5606 4850 5614
rect 4988 5676 4996 5684
rect 4972 5576 4980 5584
rect 4812 5556 4820 5564
rect 4972 5556 4980 5564
rect 4780 5496 4788 5504
rect 4972 5516 4980 5524
rect 5004 5656 5012 5664
rect 5036 5756 5044 5764
rect 5452 5756 5460 5764
rect 5548 5756 5556 5764
rect 5612 5756 5620 5764
rect 5836 5756 5844 5764
rect 5884 5756 5892 5764
rect 5084 5736 5092 5744
rect 5180 5736 5188 5744
rect 5244 5736 5252 5744
rect 5484 5736 5492 5744
rect 5068 5716 5076 5724
rect 5052 5656 5060 5664
rect 5020 5536 5028 5544
rect 5052 5536 5060 5544
rect 4828 5496 4836 5504
rect 4796 5476 4804 5484
rect 4892 5456 4900 5464
rect 4940 5496 4948 5504
rect 4972 5416 4980 5424
rect 4924 5376 4932 5384
rect 4732 5336 4740 5344
rect 4428 5316 4436 5324
rect 4492 5318 4500 5324
rect 4492 5316 4500 5318
rect 4556 5316 4564 5324
rect 4636 5316 4644 5324
rect 4380 5296 4388 5304
rect 4444 5236 4452 5244
rect 4140 5116 4148 5124
rect 4204 5116 4212 5124
rect 4076 5096 4084 5104
rect 4604 5256 4612 5264
rect 4268 5096 4276 5104
rect 4476 5096 4484 5104
rect 4524 5096 4532 5104
rect 4140 5056 4148 5064
rect 3980 4976 3988 4984
rect 4444 5056 4452 5064
rect 4412 5036 4420 5044
rect 4124 4956 4132 4964
rect 4156 4956 4164 4964
rect 3980 4918 3988 4924
rect 3980 4916 3988 4918
rect 4252 4916 4260 4924
rect 4140 4876 4148 4884
rect 3948 4816 3956 4824
rect 4108 4816 4116 4824
rect 4108 4736 4116 4744
rect 3932 4716 3940 4724
rect 3996 4716 4004 4724
rect 3980 4696 3988 4704
rect 4012 4696 4020 4704
rect 3852 4556 3860 4564
rect 3772 4536 3780 4544
rect 3852 4536 3860 4544
rect 3660 4516 3668 4524
rect 3676 4496 3684 4504
rect 3612 4296 3620 4304
rect 3788 4496 3796 4504
rect 3804 4496 3812 4504
rect 3820 4476 3828 4484
rect 3900 4656 3908 4664
rect 3916 4636 3924 4644
rect 3916 4596 3924 4604
rect 3900 4576 3908 4584
rect 3916 4536 3924 4544
rect 3868 4436 3876 4444
rect 3628 4276 3636 4284
rect 3788 4276 3796 4284
rect 3612 4236 3620 4244
rect 3724 4236 3732 4244
rect 3756 4236 3764 4244
rect 3804 4236 3812 4244
rect 3564 4196 3572 4204
rect 3500 4136 3508 4144
rect 3484 4116 3492 4124
rect 3388 3996 3396 4004
rect 3212 3876 3220 3884
rect 3340 3856 3348 3864
rect 3244 3836 3252 3844
rect 3276 3836 3284 3844
rect 2908 3736 2916 3744
rect 2892 3676 2900 3684
rect 2764 3636 2772 3644
rect 2796 3636 2804 3644
rect 2620 3576 2628 3584
rect 2492 3556 2500 3564
rect 2604 3556 2612 3564
rect 2476 3516 2484 3524
rect 2300 3476 2308 3484
rect 2444 3476 2452 3484
rect 2092 3456 2100 3464
rect 1868 3336 1876 3344
rect 2012 3416 2020 3424
rect 1948 3396 1956 3404
rect 1932 3376 1940 3384
rect 1900 3356 1908 3364
rect 2220 3456 2228 3464
rect 2588 3536 2596 3544
rect 2556 3516 2564 3524
rect 2540 3496 2548 3504
rect 2652 3536 2660 3544
rect 2620 3516 2628 3524
rect 2668 3496 2676 3504
rect 2716 3496 2724 3504
rect 2556 3476 2564 3484
rect 2604 3476 2612 3484
rect 2796 3576 2804 3584
rect 2908 3576 2916 3584
rect 2892 3536 2900 3544
rect 2860 3516 2868 3524
rect 2988 3736 2996 3744
rect 3196 3736 3204 3744
rect 2988 3716 2996 3724
rect 3052 3718 3060 3724
rect 3052 3716 3060 3718
rect 2956 3676 2964 3684
rect 3196 3676 3204 3684
rect 3036 3636 3044 3644
rect 3052 3576 3060 3584
rect 3196 3576 3204 3584
rect 2924 3556 2932 3564
rect 2940 3556 2948 3564
rect 2924 3536 2932 3544
rect 2972 3536 2980 3544
rect 2988 3536 2996 3544
rect 3278 3806 3286 3814
rect 3292 3806 3300 3814
rect 3306 3806 3314 3814
rect 3404 3976 3412 3984
rect 3468 3996 3476 4004
rect 3532 4096 3540 4104
rect 3532 4016 3540 4024
rect 3500 3976 3508 3984
rect 3548 3976 3556 3984
rect 3452 3896 3460 3904
rect 3484 3896 3492 3904
rect 3516 3896 3524 3904
rect 3532 3896 3540 3904
rect 3436 3876 3444 3884
rect 3452 3856 3460 3864
rect 3420 3816 3428 3824
rect 3372 3776 3380 3784
rect 3276 3736 3284 3744
rect 3340 3716 3348 3724
rect 3356 3716 3364 3724
rect 3004 3516 3012 3524
rect 3212 3516 3220 3524
rect 2892 3476 2900 3484
rect 3020 3476 3028 3484
rect 3132 3476 3140 3484
rect 2476 3456 2484 3464
rect 2748 3456 2756 3464
rect 3004 3456 3012 3464
rect 2668 3436 2676 3444
rect 2764 3436 2772 3444
rect 2748 3416 2756 3424
rect 2428 3396 2436 3404
rect 2172 3376 2180 3384
rect 2476 3376 2484 3384
rect 2748 3376 2756 3384
rect 2044 3336 2052 3344
rect 2140 3336 2148 3344
rect 2204 3336 2212 3344
rect 2444 3336 2452 3344
rect 1884 3256 1892 3264
rect 1884 3216 1892 3224
rect 1740 3116 1748 3124
rect 1836 3116 1844 3124
rect 1756 3096 1764 3104
rect 1820 3096 1828 3104
rect 1724 3076 1732 3084
rect 2252 3296 2260 3304
rect 2012 3256 2020 3264
rect 2012 3236 2020 3244
rect 2108 3236 2116 3244
rect 1996 3116 2004 3124
rect 1964 3096 1972 3104
rect 1980 3096 1988 3104
rect 1884 3076 1892 3084
rect 1916 3076 1924 3084
rect 1980 3076 1988 3084
rect 1708 2996 1716 3004
rect 1724 2976 1732 2984
rect 1692 2956 1700 2964
rect 1356 2936 1364 2944
rect 1580 2936 1588 2944
rect 1644 2936 1652 2944
rect 1708 2936 1716 2944
rect 1436 2916 1444 2924
rect 1628 2916 1636 2924
rect 1660 2916 1668 2924
rect 1548 2876 1556 2884
rect 1612 2876 1620 2884
rect 1548 2836 1556 2844
rect 1452 2756 1460 2764
rect 1436 2736 1444 2744
rect 1308 2696 1316 2704
rect 1132 2676 1140 2684
rect 1292 2576 1300 2584
rect 1308 2576 1316 2584
rect 1228 2536 1236 2544
rect 1132 2496 1140 2504
rect 956 2436 964 2444
rect 1036 2436 1044 2444
rect 972 2316 980 2324
rect 1052 2316 1060 2324
rect 1116 2356 1124 2364
rect 1116 2316 1124 2324
rect 1148 2476 1156 2484
rect 1260 2516 1268 2524
rect 1228 2496 1236 2504
rect 1260 2496 1268 2504
rect 1276 2456 1284 2464
rect 1180 2396 1188 2404
rect 1164 2376 1172 2384
rect 1052 2296 1060 2304
rect 1100 2296 1108 2304
rect 1132 2296 1140 2304
rect 1132 2276 1140 2284
rect 748 2196 756 2204
rect 716 2156 724 2164
rect 732 2136 740 2144
rect 1004 2256 1012 2264
rect 1260 2336 1268 2344
rect 1180 2316 1188 2324
rect 1228 2316 1236 2324
rect 1212 2276 1220 2284
rect 1148 2156 1156 2164
rect 1180 2156 1188 2164
rect 1148 2136 1156 2144
rect 668 2116 676 2124
rect 684 2116 692 2124
rect 812 2118 820 2124
rect 812 2116 820 2118
rect 1020 2116 1028 2124
rect 284 2076 292 2084
rect 620 2076 628 2084
rect 668 2076 676 2084
rect 348 1936 356 1944
rect 1244 2216 1252 2224
rect 1244 2136 1252 2144
rect 1212 2116 1220 2124
rect 1308 2296 1316 2304
rect 1420 2716 1428 2724
rect 1388 2576 1396 2584
rect 1340 2556 1348 2564
rect 1580 2716 1588 2724
rect 1612 2716 1620 2724
rect 1644 2716 1652 2724
rect 1628 2696 1636 2704
rect 1564 2676 1572 2684
rect 1500 2596 1508 2604
rect 1516 2576 1524 2584
rect 1484 2556 1492 2564
rect 1356 2516 1364 2524
rect 1340 2496 1348 2504
rect 1468 2496 1476 2504
rect 1676 2676 1684 2684
rect 1612 2616 1620 2624
rect 1612 2596 1620 2604
rect 1596 2576 1604 2584
rect 1628 2576 1636 2584
rect 1660 2576 1668 2584
rect 1628 2536 1636 2544
rect 1548 2516 1556 2524
rect 1692 2656 1700 2664
rect 1932 3056 1940 3064
rect 1836 2976 1844 2984
rect 1740 2916 1748 2924
rect 1756 2916 1764 2924
rect 1932 2940 1940 2944
rect 1852 2896 1860 2904
rect 1804 2876 1812 2884
rect 1742 2806 1750 2814
rect 1756 2806 1764 2814
rect 1770 2806 1778 2814
rect 1852 2776 1860 2784
rect 1820 2696 1828 2704
rect 1836 2696 1844 2704
rect 1788 2656 1796 2664
rect 1820 2616 1828 2624
rect 1772 2596 1780 2604
rect 1772 2556 1780 2564
rect 1788 2556 1796 2564
rect 1692 2536 1700 2544
rect 1516 2496 1524 2504
rect 1612 2496 1620 2504
rect 1484 2476 1492 2484
rect 1516 2476 1524 2484
rect 1532 2476 1540 2484
rect 1484 2396 1492 2404
rect 1340 2376 1348 2384
rect 1420 2376 1428 2384
rect 1468 2336 1476 2344
rect 1388 2316 1396 2324
rect 1372 2296 1380 2304
rect 1436 2296 1444 2304
rect 1356 2276 1364 2284
rect 1340 2236 1348 2244
rect 1324 2176 1332 2184
rect 1292 2156 1300 2164
rect 1276 2136 1284 2144
rect 1308 2136 1316 2144
rect 940 2076 948 2084
rect 1068 2076 1076 2084
rect 908 1976 916 1984
rect 652 1956 660 1964
rect 844 1956 852 1964
rect 636 1936 644 1944
rect 380 1896 388 1904
rect 428 1896 436 1904
rect 92 1856 100 1864
rect 28 1676 36 1684
rect 60 1696 68 1704
rect 12 1476 20 1484
rect 92 1536 100 1544
rect 172 1696 180 1704
rect 124 1676 132 1684
rect 140 1516 148 1524
rect 364 1876 372 1884
rect 492 1876 500 1884
rect 300 1856 308 1864
rect 460 1856 468 1864
rect 236 1756 244 1764
rect 588 1796 596 1804
rect 428 1776 436 1784
rect 524 1776 532 1784
rect 668 1936 676 1944
rect 716 1936 724 1944
rect 1020 1936 1028 1944
rect 796 1916 804 1924
rect 668 1896 676 1904
rect 636 1796 644 1804
rect 620 1776 628 1784
rect 332 1756 340 1764
rect 540 1756 548 1764
rect 220 1556 228 1564
rect 284 1556 292 1564
rect 236 1516 244 1524
rect 156 1496 164 1504
rect 220 1496 228 1504
rect 76 1476 84 1484
rect 108 1476 116 1484
rect 156 1476 164 1484
rect 268 1476 276 1484
rect 28 1456 36 1464
rect 124 1456 132 1464
rect 124 1356 132 1364
rect 12 1336 20 1344
rect 44 1316 52 1324
rect 140 1316 148 1324
rect 172 1316 180 1324
rect 236 1318 244 1324
rect 236 1316 244 1318
rect 172 1276 180 1284
rect 332 1716 340 1724
rect 444 1716 452 1724
rect 428 1636 436 1644
rect 396 1556 404 1564
rect 316 1536 324 1544
rect 412 1516 420 1524
rect 332 1496 340 1504
rect 348 1476 356 1484
rect 380 1476 388 1484
rect 300 1276 308 1284
rect 268 1256 276 1264
rect 460 1636 468 1644
rect 412 1476 420 1484
rect 540 1676 548 1684
rect 604 1676 612 1684
rect 492 1496 500 1504
rect 524 1496 532 1504
rect 540 1476 548 1484
rect 572 1496 580 1504
rect 524 1456 532 1464
rect 556 1456 564 1464
rect 476 1436 484 1444
rect 380 1356 388 1364
rect 396 1356 404 1364
rect 412 1336 420 1344
rect 460 1356 468 1364
rect 380 1316 388 1324
rect 428 1316 436 1324
rect 556 1436 564 1444
rect 540 1376 548 1384
rect 460 1316 468 1324
rect 492 1316 500 1324
rect 364 1296 372 1304
rect 444 1296 452 1304
rect 364 1256 372 1264
rect 364 1156 372 1164
rect 348 1116 356 1124
rect 492 1256 500 1264
rect 428 1116 436 1124
rect 396 1096 404 1104
rect 204 1036 212 1044
rect 220 1036 228 1044
rect 108 976 116 984
rect 44 956 52 964
rect 140 936 148 944
rect 188 936 196 944
rect 28 916 36 924
rect 92 916 100 924
rect 156 916 164 924
rect 204 916 212 924
rect 12 876 20 884
rect 60 896 68 904
rect 172 896 180 904
rect 204 896 212 904
rect 140 876 148 884
rect 76 856 84 864
rect 28 736 36 744
rect 12 696 20 704
rect 124 756 132 764
rect 76 696 84 704
rect 236 976 244 984
rect 316 1036 324 1044
rect 300 956 308 964
rect 412 996 420 1004
rect 364 936 372 944
rect 268 916 276 924
rect 412 916 420 924
rect 284 876 292 884
rect 236 776 244 784
rect 252 736 260 744
rect 284 736 292 744
rect 220 716 228 724
rect 12 596 20 604
rect 60 596 68 604
rect 172 696 180 704
rect 316 876 324 884
rect 348 876 356 884
rect 428 896 436 904
rect 396 876 404 884
rect 364 856 372 864
rect 364 776 372 784
rect 316 716 324 724
rect 300 696 308 704
rect 332 696 340 704
rect 172 676 180 684
rect 220 676 228 684
rect 252 676 260 684
rect 348 676 356 684
rect 172 576 180 584
rect 284 556 292 564
rect 140 536 148 544
rect 204 536 212 544
rect 252 536 260 544
rect 140 302 148 304
rect 140 296 148 302
rect 396 776 404 784
rect 508 1016 516 1024
rect 636 1756 644 1764
rect 764 1896 772 1904
rect 844 1916 852 1924
rect 716 1776 724 1784
rect 732 1756 740 1764
rect 780 1756 788 1764
rect 700 1736 708 1744
rect 684 1696 692 1704
rect 908 1916 916 1924
rect 1004 1916 1012 1924
rect 892 1896 900 1904
rect 908 1896 916 1904
rect 972 1896 980 1904
rect 860 1836 868 1844
rect 908 1836 916 1844
rect 892 1816 900 1824
rect 828 1776 836 1784
rect 940 1816 948 1824
rect 908 1756 916 1764
rect 924 1756 932 1764
rect 796 1736 804 1744
rect 764 1716 772 1724
rect 796 1716 804 1724
rect 892 1716 900 1724
rect 908 1596 916 1604
rect 732 1496 740 1504
rect 764 1502 772 1504
rect 764 1496 772 1502
rect 828 1496 836 1504
rect 684 1480 692 1484
rect 684 1476 692 1480
rect 572 1336 580 1344
rect 588 1336 596 1344
rect 572 1316 580 1324
rect 556 1296 564 1304
rect 572 1276 580 1284
rect 636 1336 644 1344
rect 620 1296 628 1304
rect 588 1016 596 1024
rect 604 996 612 1004
rect 556 976 564 984
rect 460 716 468 724
rect 428 696 436 704
rect 460 702 468 704
rect 460 696 468 702
rect 492 676 500 684
rect 380 596 388 604
rect 364 556 372 564
rect 588 896 596 904
rect 892 1396 900 1404
rect 684 1376 692 1384
rect 796 1316 804 1324
rect 876 1316 884 1324
rect 860 1196 868 1204
rect 1292 2056 1300 2064
rect 1228 1976 1236 1984
rect 1308 1976 1316 1984
rect 1084 1916 1092 1924
rect 1164 1916 1172 1924
rect 1212 1916 1220 1924
rect 1068 1896 1076 1904
rect 1116 1896 1124 1904
rect 1180 1896 1188 1904
rect 1036 1876 1044 1884
rect 988 1836 996 1844
rect 1052 1756 1060 1764
rect 1084 1836 1092 1844
rect 940 1736 948 1744
rect 956 1736 964 1744
rect 1068 1736 1076 1744
rect 1004 1716 1012 1724
rect 956 1696 964 1704
rect 972 1496 980 1504
rect 924 1396 932 1404
rect 1196 1876 1204 1884
rect 1244 1936 1252 1944
rect 1436 2276 1444 2284
rect 1404 2236 1412 2244
rect 1420 2196 1428 2204
rect 1660 2456 1668 2464
rect 1548 2356 1556 2364
rect 1564 2356 1572 2364
rect 1532 2316 1540 2324
rect 1548 2296 1556 2304
rect 1644 2256 1652 2264
rect 1724 2516 1732 2524
rect 1740 2516 1748 2524
rect 1836 2536 1844 2544
rect 1884 2756 1892 2764
rect 1884 2736 1892 2744
rect 1868 2616 1876 2624
rect 1932 2936 1940 2940
rect 1948 2916 1956 2924
rect 1948 2696 1956 2704
rect 2012 3096 2020 3104
rect 2028 3076 2036 3084
rect 2012 2976 2020 2984
rect 2044 2956 2052 2964
rect 2028 2936 2036 2944
rect 2028 2916 2036 2924
rect 2012 2896 2020 2904
rect 2364 3236 2372 3244
rect 2300 3136 2308 3144
rect 2188 3116 2196 3124
rect 2364 3116 2372 3124
rect 2172 3076 2180 3084
rect 2316 3076 2324 3084
rect 2092 2956 2100 2964
rect 2428 3296 2436 3304
rect 2508 3356 2516 3364
rect 2588 3356 2596 3364
rect 2636 3356 2644 3364
rect 2700 3356 2708 3364
rect 2492 3336 2500 3344
rect 2540 3336 2548 3344
rect 2604 3336 2612 3344
rect 2540 3296 2548 3304
rect 2460 3276 2468 3284
rect 2492 3276 2500 3284
rect 2412 3156 2420 3164
rect 2476 3156 2484 3164
rect 2556 3156 2564 3164
rect 2412 3136 2420 3144
rect 2444 3116 2452 3124
rect 2508 3116 2516 3124
rect 2492 3096 2500 3104
rect 2412 3076 2420 3084
rect 2460 3076 2468 3084
rect 2332 2976 2340 2984
rect 2380 2976 2388 2984
rect 2220 2956 2228 2964
rect 2300 2936 2308 2944
rect 2348 2936 2356 2944
rect 2396 2936 2404 2944
rect 2572 3096 2580 3104
rect 2572 3076 2580 3084
rect 2588 3056 2596 3064
rect 2684 3336 2692 3344
rect 2796 3376 2804 3384
rect 2764 3356 2772 3364
rect 2652 3296 2660 3304
rect 2748 3296 2756 3304
rect 2668 3276 2676 3284
rect 2620 3236 2628 3244
rect 2652 3116 2660 3124
rect 2652 3096 2660 3104
rect 2620 3076 2628 3084
rect 2604 3036 2612 3044
rect 2460 2976 2468 2984
rect 2492 2976 2500 2984
rect 2572 2976 2580 2984
rect 2444 2936 2452 2944
rect 2492 2956 2500 2964
rect 2620 2956 2628 2964
rect 2556 2936 2564 2944
rect 2588 2936 2596 2944
rect 2652 3056 2660 3064
rect 2652 3036 2660 3044
rect 2156 2918 2164 2924
rect 2156 2916 2164 2918
rect 2508 2916 2516 2924
rect 2572 2916 2580 2924
rect 2380 2896 2388 2904
rect 2524 2876 2532 2884
rect 2140 2776 2148 2784
rect 2076 2736 2084 2744
rect 2108 2736 2116 2744
rect 2044 2716 2052 2724
rect 2060 2696 2068 2704
rect 2012 2676 2020 2684
rect 1948 2656 1956 2664
rect 1980 2656 1988 2664
rect 1996 2656 2004 2664
rect 2060 2656 2068 2664
rect 1932 2556 1940 2564
rect 1884 2536 1892 2544
rect 1964 2576 1972 2584
rect 1980 2576 1988 2584
rect 2028 2576 2036 2584
rect 2076 2616 2084 2624
rect 2060 2556 2068 2564
rect 2076 2536 2084 2544
rect 1852 2516 1860 2524
rect 1916 2516 1924 2524
rect 1980 2516 1988 2524
rect 1692 2476 1700 2484
rect 1788 2476 1796 2484
rect 1836 2476 1844 2484
rect 1900 2476 1908 2484
rect 1884 2456 1892 2464
rect 1742 2406 1750 2414
rect 1756 2406 1764 2414
rect 1770 2406 1778 2414
rect 2060 2376 2068 2384
rect 2028 2356 2036 2364
rect 1900 2316 1908 2324
rect 1692 2296 1700 2304
rect 1868 2296 1876 2304
rect 1900 2296 1908 2304
rect 1948 2296 1956 2304
rect 2060 2296 2068 2304
rect 1964 2276 1972 2284
rect 2172 2696 2180 2704
rect 2124 2676 2132 2684
rect 2236 2676 2244 2684
rect 2124 2616 2132 2624
rect 2252 2596 2260 2604
rect 2140 2576 2148 2584
rect 2124 2536 2132 2544
rect 2108 2496 2116 2504
rect 2108 2276 2116 2284
rect 1868 2256 1876 2264
rect 2092 2256 2100 2264
rect 1676 2196 1684 2204
rect 1612 2156 1620 2164
rect 1660 2156 1668 2164
rect 1788 2156 1796 2164
rect 1580 2136 1588 2144
rect 1708 2136 1716 2144
rect 1676 2116 1684 2124
rect 1388 2076 1396 2084
rect 1340 2036 1348 2044
rect 1244 1916 1252 1924
rect 1324 1916 1332 1924
rect 1356 1996 1364 2004
rect 1292 1856 1300 1864
rect 1308 1776 1316 1784
rect 1228 1736 1236 1744
rect 1260 1718 1268 1724
rect 1260 1716 1268 1718
rect 1324 1716 1332 1724
rect 1116 1696 1124 1704
rect 1324 1696 1332 1704
rect 1052 1676 1060 1684
rect 1324 1656 1332 1664
rect 1068 1576 1076 1584
rect 1164 1576 1172 1584
rect 1020 1516 1028 1524
rect 1100 1556 1108 1564
rect 1052 1496 1060 1504
rect 1132 1536 1140 1544
rect 1228 1536 1236 1544
rect 1164 1516 1172 1524
rect 1148 1496 1156 1504
rect 1196 1496 1204 1504
rect 1228 1496 1236 1504
rect 1260 1496 1268 1504
rect 1148 1476 1156 1484
rect 1212 1476 1220 1484
rect 1228 1476 1236 1484
rect 1164 1456 1172 1464
rect 1148 1396 1156 1404
rect 1020 1356 1028 1364
rect 1100 1356 1108 1364
rect 1276 1436 1284 1444
rect 1180 1376 1188 1384
rect 1164 1356 1172 1364
rect 1308 1436 1316 1444
rect 1404 1956 1412 1964
rect 1372 1896 1380 1904
rect 1452 1956 1460 1964
rect 1356 1876 1364 1884
rect 1436 1876 1444 1884
rect 1356 1856 1364 1864
rect 1340 1556 1348 1564
rect 1340 1536 1348 1544
rect 1420 1836 1428 1844
rect 1372 1756 1380 1764
rect 1468 1916 1476 1924
rect 1484 1856 1492 1864
rect 1436 1756 1444 1764
rect 1452 1696 1460 1704
rect 1388 1676 1396 1684
rect 1548 2076 1556 2084
rect 1532 1736 1540 1744
rect 1500 1656 1508 1664
rect 1468 1636 1476 1644
rect 1500 1636 1508 1644
rect 1468 1516 1476 1524
rect 1404 1496 1412 1504
rect 1436 1496 1444 1504
rect 1356 1476 1364 1484
rect 1340 1456 1348 1464
rect 1420 1456 1428 1464
rect 1340 1396 1348 1404
rect 1292 1376 1300 1384
rect 1324 1356 1332 1364
rect 1132 1336 1140 1344
rect 1196 1336 1204 1344
rect 1340 1336 1348 1344
rect 908 1156 916 1164
rect 764 1136 772 1144
rect 860 1136 868 1144
rect 668 1116 676 1124
rect 732 1116 740 1124
rect 908 1116 916 1124
rect 988 1116 996 1124
rect 716 1096 724 1104
rect 860 1096 868 1104
rect 972 1096 980 1104
rect 652 1076 660 1084
rect 652 1056 660 1064
rect 748 1076 756 1084
rect 780 1076 788 1084
rect 796 1076 804 1084
rect 844 1076 852 1084
rect 876 1076 884 1084
rect 940 1076 948 1084
rect 700 1036 708 1044
rect 748 1016 756 1024
rect 764 1016 772 1024
rect 668 976 676 984
rect 652 936 660 944
rect 812 1036 820 1044
rect 828 1016 836 1024
rect 844 936 852 944
rect 956 1016 964 1024
rect 940 956 948 964
rect 988 1016 996 1024
rect 1484 1476 1492 1484
rect 1596 1956 1604 1964
rect 1596 1936 1604 1944
rect 1804 2096 1812 2104
rect 1742 2006 1750 2014
rect 1756 2006 1764 2014
rect 1770 2006 1778 2014
rect 1740 1896 1748 1904
rect 1788 1896 1796 1904
rect 1852 2156 1860 2164
rect 1852 2116 1860 2124
rect 1900 2236 1908 2244
rect 2092 2236 2100 2244
rect 2108 2136 2116 2144
rect 1932 2116 1940 2124
rect 1884 2096 1892 2104
rect 1948 2096 1956 2104
rect 1868 2076 1876 2084
rect 1820 2036 1828 2044
rect 1676 1876 1684 1884
rect 1772 1876 1780 1884
rect 1836 1836 1844 1844
rect 1660 1756 1668 1764
rect 1692 1756 1700 1764
rect 1836 1796 1844 1804
rect 2460 2796 2468 2804
rect 2300 2776 2308 2784
rect 2364 2716 2372 2724
rect 2412 2676 2420 2684
rect 2380 2656 2388 2664
rect 2316 2636 2324 2644
rect 2220 2536 2228 2544
rect 2284 2536 2292 2544
rect 2252 2516 2260 2524
rect 2236 2316 2244 2324
rect 2252 2296 2260 2304
rect 2172 2176 2180 2184
rect 2156 2156 2164 2164
rect 2172 2156 2180 2164
rect 2268 2216 2276 2224
rect 2188 2136 2196 2144
rect 2172 2116 2180 2124
rect 2140 1936 2148 1944
rect 1948 1896 1956 1904
rect 1932 1876 1940 1884
rect 2044 1876 2052 1884
rect 1868 1776 1876 1784
rect 1836 1756 1844 1764
rect 1964 1756 1972 1764
rect 1692 1736 1700 1744
rect 1820 1736 1828 1744
rect 1724 1716 1732 1724
rect 1708 1696 1716 1704
rect 1596 1676 1604 1684
rect 1644 1676 1652 1684
rect 1548 1596 1556 1604
rect 1676 1616 1684 1624
rect 1742 1606 1750 1614
rect 1756 1606 1764 1614
rect 1770 1606 1778 1614
rect 1692 1556 1700 1564
rect 1708 1556 1716 1564
rect 1548 1536 1556 1544
rect 1580 1536 1588 1544
rect 1516 1496 1524 1504
rect 1564 1496 1572 1504
rect 1580 1456 1588 1464
rect 1596 1456 1604 1464
rect 1500 1436 1508 1444
rect 1532 1436 1540 1444
rect 1484 1396 1492 1404
rect 1468 1376 1476 1384
rect 1484 1336 1492 1344
rect 1372 1316 1380 1324
rect 1676 1516 1684 1524
rect 1836 1576 1844 1584
rect 1900 1718 1908 1724
rect 1900 1716 1908 1718
rect 2028 1716 2036 1724
rect 2012 1636 2020 1644
rect 1708 1516 1716 1524
rect 1756 1516 1764 1524
rect 1804 1516 1812 1524
rect 1772 1496 1780 1504
rect 1708 1476 1716 1484
rect 1820 1476 1828 1484
rect 1612 1376 1620 1384
rect 1596 1336 1604 1344
rect 1708 1416 1716 1424
rect 1692 1376 1700 1384
rect 1612 1316 1620 1324
rect 1052 1296 1060 1304
rect 1276 1296 1284 1304
rect 1404 1296 1412 1304
rect 1436 1296 1444 1304
rect 1596 1296 1604 1304
rect 1660 1296 1668 1304
rect 1020 1196 1028 1204
rect 1020 1136 1028 1144
rect 1036 1076 1044 1084
rect 780 916 788 924
rect 876 916 884 924
rect 908 916 916 924
rect 684 896 692 904
rect 636 876 644 884
rect 796 876 804 884
rect 860 876 868 884
rect 972 876 980 884
rect 620 856 628 864
rect 588 776 596 784
rect 524 756 532 764
rect 684 716 692 724
rect 908 696 916 704
rect 700 676 708 684
rect 620 656 628 664
rect 476 636 484 644
rect 508 636 516 644
rect 396 576 404 584
rect 428 556 436 564
rect 444 536 452 544
rect 348 516 356 524
rect 524 516 532 524
rect 252 496 260 504
rect 332 496 340 504
rect 412 496 420 504
rect 492 496 500 504
rect 524 496 532 504
rect 236 336 244 344
rect 204 296 212 304
rect 812 656 820 664
rect 700 516 708 524
rect 780 516 788 524
rect 636 496 644 504
rect 572 436 580 444
rect 764 436 772 444
rect 348 336 356 344
rect 364 336 372 344
rect 252 316 260 324
rect 316 316 324 324
rect 92 256 100 264
rect 12 216 20 224
rect 252 276 260 284
rect 28 156 36 164
rect 76 156 84 164
rect 140 156 148 164
rect 60 136 68 144
rect 268 256 276 264
rect 316 256 324 264
rect 156 136 164 144
rect 316 136 324 144
rect 348 296 356 304
rect 348 156 356 164
rect 76 116 84 124
rect 188 96 196 104
rect 236 96 244 104
rect 300 96 308 104
rect 444 316 452 324
rect 572 336 580 344
rect 620 336 628 344
rect 764 336 772 344
rect 492 316 500 324
rect 396 296 404 304
rect 444 296 452 304
rect 396 276 404 284
rect 396 196 404 204
rect 588 316 596 324
rect 540 296 548 304
rect 716 302 724 304
rect 716 296 724 302
rect 460 156 468 164
rect 508 276 516 284
rect 524 256 532 264
rect 620 256 628 264
rect 652 256 660 264
rect 588 176 596 184
rect 588 136 596 144
rect 716 216 724 224
rect 716 156 724 164
rect 620 136 628 144
rect 428 116 436 124
rect 476 116 484 124
rect 604 116 612 124
rect 668 116 676 124
rect 732 116 740 124
rect 1020 956 1028 964
rect 1100 1136 1108 1144
rect 1084 1056 1092 1064
rect 1036 936 1044 944
rect 1004 896 1012 904
rect 1164 1076 1172 1084
rect 1212 1076 1220 1084
rect 1196 1056 1204 1064
rect 1116 1016 1124 1024
rect 1100 896 1108 904
rect 1468 1276 1476 1284
rect 1564 1276 1572 1284
rect 1276 1176 1284 1184
rect 1276 1136 1284 1144
rect 1228 1036 1236 1044
rect 1164 916 1172 924
rect 1660 1176 1668 1184
rect 1580 1156 1588 1164
rect 1724 1276 1732 1284
rect 1742 1206 1750 1214
rect 1756 1206 1764 1214
rect 1770 1206 1778 1214
rect 1948 1556 1956 1564
rect 1868 1536 1876 1544
rect 1916 1536 1924 1544
rect 1884 1496 1892 1504
rect 1900 1456 1908 1464
rect 1948 1456 1956 1464
rect 2060 1836 2068 1844
rect 2124 1836 2132 1844
rect 2060 1796 2068 1804
rect 2044 1496 2052 1504
rect 2092 1736 2100 1744
rect 2076 1716 2084 1724
rect 2076 1696 2084 1704
rect 2092 1676 2100 1684
rect 2076 1496 2084 1504
rect 1964 1376 1972 1384
rect 1852 1318 1860 1324
rect 1852 1316 1860 1318
rect 1916 1316 1924 1324
rect 1948 1316 1956 1324
rect 1916 1296 1924 1304
rect 1980 1296 1988 1304
rect 1980 1276 1988 1284
rect 1932 1156 1940 1164
rect 1548 1116 1556 1124
rect 1756 1116 1764 1124
rect 1324 1096 1332 1104
rect 1452 1096 1460 1104
rect 1356 1076 1364 1084
rect 1436 1076 1444 1084
rect 1340 1056 1348 1064
rect 1388 1056 1396 1064
rect 1484 1076 1492 1084
rect 1564 1076 1572 1084
rect 1660 1076 1668 1084
rect 1708 1076 1716 1084
rect 1500 1056 1508 1064
rect 1404 1036 1412 1044
rect 1452 1036 1460 1044
rect 1292 1016 1300 1024
rect 1308 996 1316 1004
rect 1260 976 1268 984
rect 1244 936 1252 944
rect 1276 936 1284 944
rect 1484 1016 1492 1024
rect 1420 996 1428 1004
rect 1468 996 1476 1004
rect 1532 996 1540 1004
rect 1484 976 1492 984
rect 1452 956 1460 964
rect 1388 936 1396 944
rect 1420 936 1428 944
rect 1212 916 1220 924
rect 1228 916 1236 924
rect 1292 916 1300 924
rect 1340 916 1348 924
rect 1388 916 1396 924
rect 1180 896 1188 904
rect 1212 896 1220 904
rect 1260 896 1268 904
rect 1356 896 1364 904
rect 1228 856 1236 864
rect 1292 736 1300 744
rect 1036 696 1044 704
rect 1436 916 1444 924
rect 1340 716 1348 724
rect 1372 716 1380 724
rect 1388 696 1396 704
rect 1196 676 1204 684
rect 1228 676 1236 684
rect 1500 956 1508 964
rect 1596 956 1604 964
rect 1612 936 1620 944
rect 1628 936 1636 944
rect 1548 896 1556 904
rect 1660 916 1668 924
rect 1452 876 1460 884
rect 1644 876 1652 884
rect 1500 756 1508 764
rect 1580 756 1588 764
rect 1532 716 1540 724
rect 1644 716 1652 724
rect 1436 696 1444 704
rect 1452 680 1460 684
rect 1452 676 1460 680
rect 1500 676 1508 684
rect 924 596 932 604
rect 988 596 996 604
rect 1484 656 1492 664
rect 1260 636 1268 644
rect 1292 636 1300 644
rect 1148 556 1156 564
rect 1132 536 1140 544
rect 844 516 852 524
rect 812 496 820 504
rect 812 436 820 444
rect 844 236 852 244
rect 876 296 884 304
rect 1004 302 1012 304
rect 1004 296 1012 302
rect 876 236 884 244
rect 860 216 868 224
rect 844 176 852 184
rect 812 136 820 144
rect 828 136 836 144
rect 796 116 804 124
rect 1244 576 1252 584
rect 1404 576 1412 584
rect 1708 976 1716 984
rect 1676 896 1684 904
rect 1724 896 1732 904
rect 1836 1056 1844 1064
rect 1756 876 1764 884
rect 1708 836 1716 844
rect 1740 836 1748 844
rect 1676 716 1684 724
rect 1742 806 1750 814
rect 1756 806 1764 814
rect 1770 806 1778 814
rect 1804 716 1812 724
rect 1548 696 1556 704
rect 1628 696 1636 704
rect 1660 696 1668 704
rect 1676 696 1684 704
rect 1772 696 1780 704
rect 1788 696 1796 704
rect 1692 656 1700 664
rect 2060 1396 2068 1404
rect 2028 1376 2036 1384
rect 2124 1416 2132 1424
rect 2268 1956 2276 1964
rect 2220 1916 2228 1924
rect 2156 1676 2164 1684
rect 2204 1896 2212 1904
rect 2188 1876 2196 1884
rect 2188 1856 2196 1864
rect 2236 1816 2244 1824
rect 2268 1756 2276 1764
rect 2204 1736 2212 1744
rect 2188 1696 2196 1704
rect 2204 1676 2212 1684
rect 2364 2536 2372 2544
rect 2348 2516 2356 2524
rect 2364 2516 2372 2524
rect 2316 2396 2324 2404
rect 2348 2236 2356 2244
rect 2316 2116 2324 2124
rect 2300 2016 2308 2024
rect 2444 2636 2452 2644
rect 2796 3296 2804 3304
rect 2844 3416 2852 3424
rect 2940 3396 2948 3404
rect 2876 3376 2884 3384
rect 2924 3336 2932 3344
rect 2956 3336 2964 3344
rect 2972 3340 2980 3344
rect 2972 3336 2980 3340
rect 2988 3336 2996 3344
rect 2876 3296 2884 3304
rect 2780 3236 2788 3244
rect 2812 3236 2820 3244
rect 2684 3156 2692 3164
rect 2908 3196 2916 3204
rect 2940 3196 2948 3204
rect 2796 3156 2804 3164
rect 2716 3096 2724 3104
rect 2764 3116 2772 3124
rect 2780 3096 2788 3104
rect 2828 3116 2836 3124
rect 2924 3076 2932 3084
rect 2892 3036 2900 3044
rect 2684 2916 2692 2924
rect 2940 2936 2948 2944
rect 2700 2896 2708 2904
rect 2924 2916 2932 2924
rect 2892 2896 2900 2904
rect 2908 2876 2916 2884
rect 2908 2856 2916 2864
rect 2876 2836 2884 2844
rect 2860 2796 2868 2804
rect 3196 3336 3204 3344
rect 3260 3656 3268 3664
rect 3436 3756 3444 3764
rect 3404 3736 3412 3744
rect 3580 3876 3588 3884
rect 3564 3856 3572 3864
rect 3596 3856 3604 3864
rect 3580 3836 3588 3844
rect 3532 3816 3540 3824
rect 3468 3756 3476 3764
rect 3468 3736 3476 3744
rect 3436 3716 3444 3724
rect 3548 3776 3556 3784
rect 3516 3736 3524 3744
rect 3564 3756 3572 3764
rect 3788 4176 3796 4184
rect 3708 4156 3716 4164
rect 3756 4156 3764 4164
rect 3836 4336 3844 4344
rect 3884 4336 3892 4344
rect 3868 4236 3876 4244
rect 3916 4156 3924 4164
rect 3964 4676 3972 4684
rect 3948 4616 3956 4624
rect 3948 4576 3956 4584
rect 3948 4516 3956 4524
rect 3996 4516 4004 4524
rect 3980 4496 3988 4504
rect 4060 4636 4068 4644
rect 4044 4576 4052 4584
rect 4028 4536 4036 4544
rect 4028 4516 4036 4524
rect 3964 4456 3972 4464
rect 3964 4436 3972 4444
rect 3948 4356 3956 4364
rect 4012 4456 4020 4464
rect 4044 4396 4052 4404
rect 4044 4376 4052 4384
rect 4012 4336 4020 4344
rect 3996 4316 4004 4324
rect 3948 4276 3956 4284
rect 3948 4236 3956 4244
rect 4012 4196 4020 4204
rect 3724 4116 3732 4124
rect 3772 4116 3780 4124
rect 3820 4116 3828 4124
rect 3948 4116 3956 4124
rect 3884 4076 3892 4084
rect 3692 4056 3700 4064
rect 3660 3996 3668 4004
rect 3628 3916 3636 3924
rect 3692 3916 3700 3924
rect 3708 3916 3716 3924
rect 3740 3916 3748 3924
rect 3756 3916 3764 3924
rect 3788 3916 3796 3924
rect 3628 3876 3636 3884
rect 3708 3896 3716 3904
rect 3724 3896 3732 3904
rect 3724 3876 3732 3884
rect 3708 3836 3716 3844
rect 3724 3776 3732 3784
rect 3772 3896 3780 3904
rect 3820 3916 3828 3924
rect 3852 3896 3860 3904
rect 3884 3896 3892 3904
rect 3788 3856 3796 3864
rect 3916 4096 3924 4104
rect 3932 4016 3940 4024
rect 3836 3836 3844 3844
rect 3900 3836 3908 3844
rect 3612 3756 3620 3764
rect 3628 3756 3636 3764
rect 3660 3756 3668 3764
rect 3676 3756 3684 3764
rect 3756 3756 3764 3764
rect 3580 3716 3588 3724
rect 3628 3716 3636 3724
rect 3644 3716 3652 3724
rect 3788 3736 3796 3744
rect 3948 3736 3956 3744
rect 3708 3716 3716 3724
rect 3916 3716 3924 3724
rect 3500 3656 3508 3664
rect 3276 3636 3284 3644
rect 3452 3636 3460 3644
rect 3580 3616 3588 3624
rect 3516 3576 3524 3584
rect 3436 3556 3444 3564
rect 3356 3536 3364 3544
rect 3388 3516 3396 3524
rect 3420 3516 3428 3524
rect 3596 3516 3604 3524
rect 3244 3496 3252 3504
rect 3356 3496 3364 3504
rect 3516 3496 3524 3504
rect 3260 3456 3268 3464
rect 3388 3456 3396 3464
rect 3340 3436 3348 3444
rect 3278 3406 3286 3414
rect 3292 3406 3300 3414
rect 3306 3406 3314 3414
rect 3468 3436 3476 3444
rect 3436 3416 3444 3424
rect 3340 3376 3348 3384
rect 3388 3376 3396 3384
rect 3372 3356 3380 3364
rect 3420 3356 3428 3364
rect 3052 3096 3060 3104
rect 3260 3316 3268 3324
rect 3116 3296 3124 3304
rect 3164 3296 3172 3304
rect 3500 3436 3508 3444
rect 3564 3436 3572 3444
rect 3500 3376 3508 3384
rect 3500 3356 3508 3364
rect 3484 3316 3492 3324
rect 3356 3296 3364 3304
rect 3340 3216 3348 3224
rect 3164 3096 3172 3104
rect 3180 3096 3188 3104
rect 3132 3076 3140 3084
rect 3020 3056 3028 3064
rect 2988 2976 2996 2984
rect 3196 3076 3204 3084
rect 3324 3136 3332 3144
rect 3564 3376 3572 3384
rect 3532 3336 3540 3344
rect 3372 3276 3380 3284
rect 3420 3276 3428 3284
rect 3532 3156 3540 3164
rect 3452 3136 3460 3144
rect 3468 3136 3476 3144
rect 3420 3116 3428 3124
rect 3500 3116 3508 3124
rect 3740 3556 3748 3564
rect 3772 3556 3780 3564
rect 3804 3556 3812 3564
rect 3852 3556 3860 3564
rect 3628 3536 3636 3544
rect 3724 3536 3732 3544
rect 3628 3476 3636 3484
rect 3660 3456 3668 3464
rect 3676 3456 3684 3464
rect 3644 3416 3652 3424
rect 3692 3416 3700 3424
rect 3708 3356 3716 3364
rect 3660 3336 3668 3344
rect 3628 3296 3636 3304
rect 3820 3516 3828 3524
rect 3884 3516 3892 3524
rect 3772 3496 3780 3504
rect 3852 3476 3860 3484
rect 3868 3476 3876 3484
rect 3740 3436 3748 3444
rect 3756 3436 3764 3444
rect 3804 3436 3812 3444
rect 3788 3376 3796 3384
rect 3804 3376 3812 3384
rect 3868 3416 3876 3424
rect 3820 3356 3828 3364
rect 3852 3356 3860 3364
rect 4092 4536 4100 4544
rect 4108 4456 4116 4464
rect 4076 4436 4084 4444
rect 4076 4396 4084 4404
rect 4060 4336 4068 4344
rect 4076 4296 4084 4304
rect 4156 4836 4164 4844
rect 4284 4776 4292 4784
rect 4156 4716 4164 4724
rect 4220 4702 4228 4704
rect 4220 4696 4228 4702
rect 4236 4596 4244 4604
rect 4220 4576 4228 4584
rect 4364 4916 4372 4924
rect 4364 4896 4372 4904
rect 4396 4836 4404 4844
rect 4348 4796 4356 4804
rect 4588 4936 4596 4944
rect 4636 5156 4644 5164
rect 4732 5136 4740 5144
rect 5020 5416 5028 5424
rect 5004 5376 5012 5384
rect 5004 5356 5012 5364
rect 4764 5336 4772 5344
rect 4988 5336 4996 5344
rect 4748 5116 4756 5124
rect 4716 5096 4724 5104
rect 4700 5076 4708 5084
rect 4748 5076 4756 5084
rect 4652 5056 4660 5064
rect 4636 5036 4644 5044
rect 4700 5056 4708 5064
rect 4748 4996 4756 5004
rect 4716 4956 4724 4964
rect 4780 5236 4788 5244
rect 4814 5206 4822 5214
rect 4828 5206 4836 5214
rect 4842 5206 4850 5214
rect 4828 5176 4836 5184
rect 4876 5156 4884 5164
rect 4796 5116 4804 5124
rect 4908 5296 4916 5304
rect 4940 5256 4948 5264
rect 4908 5176 4916 5184
rect 4892 5136 4900 5144
rect 5020 5336 5028 5344
rect 5068 5516 5076 5524
rect 5068 5496 5076 5504
rect 5132 5716 5140 5724
rect 5180 5716 5188 5724
rect 5212 5696 5220 5704
rect 5372 5696 5380 5704
rect 5500 5716 5508 5724
rect 5516 5696 5524 5704
rect 5116 5676 5124 5684
rect 5388 5676 5396 5684
rect 5100 5536 5108 5544
rect 5164 5536 5172 5544
rect 5084 5456 5092 5464
rect 5068 5416 5076 5424
rect 5484 5676 5492 5684
rect 5468 5656 5476 5664
rect 5420 5636 5428 5644
rect 5532 5636 5540 5644
rect 5388 5576 5396 5584
rect 5148 5496 5156 5504
rect 5180 5496 5188 5504
rect 5388 5496 5396 5504
rect 5132 5476 5140 5484
rect 5116 5456 5124 5464
rect 5212 5456 5220 5464
rect 5228 5456 5236 5464
rect 5148 5416 5156 5424
rect 5196 5416 5204 5424
rect 5100 5376 5108 5384
rect 5116 5376 5124 5384
rect 5196 5356 5204 5364
rect 5212 5356 5220 5364
rect 5132 5316 5140 5324
rect 5180 5316 5188 5324
rect 5052 5296 5060 5304
rect 5196 5296 5204 5304
rect 4924 5116 4932 5124
rect 5020 5116 5028 5124
rect 5036 5096 5044 5104
rect 5148 5176 5156 5184
rect 5244 5436 5252 5444
rect 5276 5456 5284 5464
rect 5228 5316 5236 5324
rect 5436 5456 5444 5464
rect 5564 5656 5572 5664
rect 5612 5736 5620 5744
rect 5612 5716 5620 5724
rect 5660 5696 5668 5704
rect 5628 5596 5636 5604
rect 5580 5576 5588 5584
rect 5692 5716 5700 5724
rect 5708 5676 5716 5684
rect 5836 5736 5844 5744
rect 5900 5736 5908 5744
rect 6092 5736 6100 5744
rect 5772 5716 5780 5724
rect 5820 5716 5828 5724
rect 5788 5696 5796 5704
rect 5804 5696 5812 5704
rect 5756 5656 5764 5664
rect 5724 5616 5732 5624
rect 5852 5696 5860 5704
rect 5868 5676 5876 5684
rect 5916 5676 5924 5684
rect 5836 5656 5844 5664
rect 5804 5636 5812 5644
rect 5884 5636 5892 5644
rect 5740 5596 5748 5604
rect 5756 5596 5764 5604
rect 5740 5576 5748 5584
rect 5772 5536 5780 5544
rect 5804 5556 5812 5564
rect 5836 5536 5844 5544
rect 5868 5516 5876 5524
rect 5788 5496 5796 5504
rect 5852 5496 5860 5504
rect 5916 5596 5924 5604
rect 5900 5556 5908 5564
rect 5900 5496 5908 5504
rect 5516 5476 5524 5484
rect 5676 5476 5684 5484
rect 5756 5476 5764 5484
rect 5580 5456 5588 5464
rect 5884 5456 5892 5464
rect 5980 5716 5988 5724
rect 5948 5636 5956 5644
rect 5996 5616 6004 5624
rect 6028 5516 6036 5524
rect 5996 5496 6004 5504
rect 6028 5496 6036 5504
rect 6204 5776 6212 5784
rect 6188 5756 6196 5764
rect 6572 5756 6580 5764
rect 6780 5756 6788 5764
rect 7052 5756 7060 5764
rect 7324 5756 7332 5764
rect 6364 5736 6372 5744
rect 6444 5736 6452 5744
rect 6652 5736 6660 5744
rect 6908 5736 6916 5744
rect 7116 5736 7124 5744
rect 7164 5736 7172 5744
rect 7340 5736 7348 5744
rect 7612 5736 7620 5744
rect 7964 5736 7972 5744
rect 7996 5736 8004 5744
rect 6076 5716 6084 5724
rect 6316 5716 6324 5724
rect 6716 5718 6724 5724
rect 6716 5716 6724 5718
rect 6748 5716 6756 5724
rect 6092 5676 6100 5684
rect 6060 5656 6068 5664
rect 6188 5576 6196 5584
rect 6140 5516 6148 5524
rect 6204 5536 6212 5544
rect 6508 5536 6516 5544
rect 6700 5536 6708 5544
rect 6892 5536 6900 5544
rect 6588 5516 6596 5524
rect 6620 5516 6628 5524
rect 6684 5516 6692 5524
rect 6540 5496 6548 5504
rect 6572 5496 6580 5504
rect 6604 5496 6612 5504
rect 6636 5496 6644 5504
rect 6684 5496 6692 5504
rect 6044 5476 6052 5484
rect 6108 5456 6116 5464
rect 5548 5436 5556 5444
rect 5708 5436 5716 5444
rect 5932 5436 5940 5444
rect 5948 5436 5956 5444
rect 5340 5356 5348 5364
rect 5372 5356 5380 5364
rect 5292 5336 5300 5344
rect 5436 5336 5444 5344
rect 5500 5336 5508 5344
rect 5548 5336 5556 5344
rect 5564 5336 5572 5344
rect 5244 5296 5252 5304
rect 5340 5316 5348 5324
rect 5420 5316 5428 5324
rect 5436 5316 5444 5324
rect 5484 5316 5492 5324
rect 5340 5276 5348 5284
rect 5276 5176 5284 5184
rect 5404 5116 5412 5124
rect 5164 5102 5172 5104
rect 5164 5096 5172 5102
rect 5388 5096 5396 5104
rect 5420 5096 5428 5104
rect 5452 5096 5460 5104
rect 5900 5416 5908 5424
rect 6188 5416 6196 5424
rect 6044 5376 6052 5384
rect 5516 5316 5524 5324
rect 5660 5316 5668 5324
rect 5692 5316 5700 5324
rect 5772 5316 5780 5324
rect 5532 5116 5540 5124
rect 4796 5076 4804 5084
rect 4972 5076 4980 5084
rect 5100 5076 5108 5084
rect 5260 5076 5268 5084
rect 5436 5076 5444 5084
rect 5500 5076 5508 5084
rect 5516 5076 5524 5084
rect 4940 5056 4948 5064
rect 4780 5036 4788 5044
rect 4876 5036 4884 5044
rect 4780 4976 4788 4984
rect 4908 4976 4916 4984
rect 4764 4936 4772 4944
rect 4620 4896 4628 4904
rect 4604 4836 4612 4844
rect 4476 4776 4484 4784
rect 4492 4776 4500 4784
rect 4444 4756 4452 4764
rect 4476 4756 4484 4764
rect 4348 4696 4356 4704
rect 4364 4676 4372 4684
rect 4412 4676 4420 4684
rect 4492 4696 4500 4704
rect 4556 4696 4564 4704
rect 4588 4696 4596 4704
rect 4604 4696 4612 4704
rect 4460 4676 4468 4684
rect 4524 4676 4532 4684
rect 4556 4676 4564 4684
rect 4716 4876 4724 4884
rect 4748 4876 4756 4884
rect 4796 4876 4804 4884
rect 4636 4796 4644 4804
rect 4732 4716 4740 4724
rect 4814 4806 4822 4814
rect 4828 4806 4836 4814
rect 4842 4806 4850 4814
rect 5228 5056 5236 5064
rect 5308 5056 5316 5064
rect 4972 4936 4980 4944
rect 5068 4936 5076 4944
rect 5196 4916 5204 4924
rect 5132 4876 5140 4884
rect 5004 4836 5012 4844
rect 5244 4836 5252 4844
rect 4940 4816 4948 4824
rect 5148 4816 5156 4824
rect 4908 4756 4916 4764
rect 5004 4756 5012 4764
rect 5020 4756 5028 4764
rect 5052 4756 5060 4764
rect 5116 4756 5124 4764
rect 5164 4756 5172 4764
rect 4828 4716 4836 4724
rect 4684 4696 4692 4704
rect 4700 4696 4708 4704
rect 4716 4696 4724 4704
rect 4748 4696 4756 4704
rect 4684 4676 4692 4684
rect 4508 4656 4516 4664
rect 4572 4656 4580 4664
rect 4588 4656 4596 4664
rect 4652 4656 4660 4664
rect 4668 4656 4676 4664
rect 4348 4636 4356 4644
rect 4444 4636 4452 4644
rect 4412 4616 4420 4624
rect 4380 4596 4388 4604
rect 4332 4576 4340 4584
rect 4316 4556 4324 4564
rect 4252 4536 4260 4544
rect 4284 4536 4292 4544
rect 4348 4536 4356 4544
rect 4172 4516 4180 4524
rect 4188 4496 4196 4504
rect 4140 4436 4148 4444
rect 4220 4356 4228 4364
rect 4188 4296 4196 4304
rect 4268 4516 4276 4524
rect 4348 4516 4356 4524
rect 4300 4416 4308 4424
rect 4316 4336 4324 4344
rect 4284 4316 4292 4324
rect 4316 4276 4324 4284
rect 4124 4216 4132 4224
rect 4028 4176 4036 4184
rect 4156 4156 4164 4164
rect 4012 4116 4020 4124
rect 3996 4096 4004 4104
rect 3980 4016 3988 4024
rect 4076 4056 4084 4064
rect 4060 3996 4068 4004
rect 4028 3976 4036 3984
rect 4060 3896 4068 3904
rect 4076 3896 4084 3904
rect 3980 3876 3988 3884
rect 4028 3856 4036 3864
rect 4268 4196 4276 4204
rect 4348 4156 4356 4164
rect 4428 4576 4436 4584
rect 4508 4576 4516 4584
rect 4636 4636 4644 4644
rect 4588 4596 4596 4604
rect 4764 4676 4772 4684
rect 4940 4716 4948 4724
rect 4988 4716 4996 4724
rect 5036 4716 5044 4724
rect 5052 4716 5060 4724
rect 5180 4716 5188 4724
rect 5276 4716 5284 4724
rect 4748 4656 4756 4664
rect 4860 4656 4868 4664
rect 4972 4656 4980 4664
rect 5036 4656 5044 4664
rect 4764 4616 4772 4624
rect 4620 4516 4628 4524
rect 4556 4496 4564 4504
rect 4556 4476 4564 4484
rect 4460 4436 4468 4444
rect 4460 4336 4468 4344
rect 4476 4336 4484 4344
rect 4444 4316 4452 4324
rect 4396 4196 4404 4204
rect 4444 4176 4452 4184
rect 4380 4156 4388 4164
rect 4412 4156 4420 4164
rect 4300 4116 4308 4124
rect 4332 4116 4340 4124
rect 4364 4116 4372 4124
rect 4236 4096 4244 4104
rect 4204 3902 4212 3904
rect 4204 3896 4212 3902
rect 4108 3876 4116 3884
rect 4092 3816 4100 3824
rect 4012 3756 4020 3764
rect 4172 3856 4180 3864
rect 4140 3836 4148 3844
rect 4204 3816 4212 3824
rect 4204 3756 4212 3764
rect 4220 3756 4228 3764
rect 4076 3736 4084 3744
rect 3980 3636 3988 3644
rect 3964 3596 3972 3604
rect 3964 3536 3972 3544
rect 3932 3456 3940 3464
rect 3916 3376 3924 3384
rect 3900 3336 3908 3344
rect 3916 3336 3924 3344
rect 4140 3496 4148 3504
rect 4156 3496 4164 3504
rect 3996 3476 4004 3484
rect 4060 3476 4068 3484
rect 4108 3476 4116 3484
rect 4028 3456 4036 3464
rect 3996 3396 4004 3404
rect 4060 3356 4068 3364
rect 4156 3376 4164 3384
rect 4204 3376 4212 3384
rect 4012 3336 4020 3344
rect 4124 3336 4132 3344
rect 3756 3316 3764 3324
rect 3916 3316 3924 3324
rect 4172 3356 4180 3364
rect 4268 3996 4276 4004
rect 4316 4056 4324 4064
rect 4316 3996 4324 4004
rect 4348 3996 4356 4004
rect 4684 4516 4692 4524
rect 4716 4456 4724 4464
rect 4636 4436 4644 4444
rect 4588 4316 4596 4324
rect 4924 4516 4932 4524
rect 4780 4476 4788 4484
rect 4972 4476 4980 4484
rect 4876 4456 4884 4464
rect 5100 4696 5108 4704
rect 5116 4676 5124 4684
rect 5164 4676 5172 4684
rect 5084 4556 5092 4564
rect 5068 4536 5076 4544
rect 5116 4536 5124 4544
rect 5132 4516 5140 4524
rect 5052 4496 5060 4504
rect 5212 4676 5220 4684
rect 5196 4636 5204 4644
rect 5180 4536 5188 4544
rect 5068 4476 5076 4484
rect 4732 4436 4740 4444
rect 4844 4436 4852 4444
rect 4876 4436 4884 4444
rect 5004 4436 5012 4444
rect 4588 4296 4596 4304
rect 4652 4302 4660 4304
rect 4652 4296 4660 4302
rect 4700 4296 4708 4304
rect 4524 4256 4532 4264
rect 4508 4216 4516 4224
rect 4492 4196 4500 4204
rect 4492 4116 4500 4124
rect 4460 4076 4468 4084
rect 4508 4076 4516 4084
rect 4364 3956 4372 3964
rect 4476 3996 4484 4004
rect 4412 3976 4420 3984
rect 4348 3936 4356 3944
rect 4332 3896 4340 3904
rect 4332 3836 4340 3844
rect 4300 3756 4308 3764
rect 4396 3936 4404 3944
rect 4396 3796 4404 3804
rect 4428 3796 4436 3804
rect 4412 3736 4420 3744
rect 4332 3696 4340 3704
rect 4268 3636 4276 3644
rect 4300 3596 4308 3604
rect 4252 3516 4260 3524
rect 4268 3516 4276 3524
rect 4236 3336 4244 3344
rect 4204 3316 4212 3324
rect 4332 3596 4340 3604
rect 4380 3536 4388 3544
rect 4476 3876 4484 3884
rect 4556 4176 4564 4184
rect 4540 4156 4548 4164
rect 4540 4016 4548 4024
rect 4588 4076 4596 4084
rect 4572 3876 4580 3884
rect 4540 3836 4548 3844
rect 4814 4406 4822 4414
rect 4828 4406 4836 4414
rect 4842 4406 4850 4414
rect 4844 4296 4852 4304
rect 4700 4236 4708 4244
rect 4780 4236 4788 4244
rect 4860 4236 4868 4244
rect 4764 4216 4772 4224
rect 4844 4196 4852 4204
rect 4716 4156 4724 4164
rect 4796 4156 4804 4164
rect 4860 4176 4868 4184
rect 4988 4416 4996 4424
rect 4892 4316 4900 4324
rect 5132 4336 5140 4344
rect 5180 4336 5188 4344
rect 4988 4276 4996 4284
rect 5036 4276 5044 4284
rect 5148 4276 5156 4284
rect 4972 4256 4980 4264
rect 4956 4236 4964 4244
rect 4940 4216 4948 4224
rect 4924 4176 4932 4184
rect 4972 4176 4980 4184
rect 4940 4156 4948 4164
rect 4684 4136 4692 4144
rect 4700 4136 4708 4144
rect 4780 4136 4788 4144
rect 4876 4136 4884 4144
rect 4972 4136 4980 4144
rect 4684 4056 4692 4064
rect 4668 3996 4676 4004
rect 4652 3936 4660 3944
rect 4636 3836 4644 3844
rect 4684 3836 4692 3844
rect 4556 3796 4564 3804
rect 4620 3796 4628 3804
rect 4540 3776 4548 3784
rect 4652 3756 4660 3764
rect 4620 3736 4628 3744
rect 4748 4076 4756 4084
rect 4748 3996 4756 4004
rect 4732 3956 4740 3964
rect 4700 3776 4708 3784
rect 4716 3756 4724 3764
rect 4876 4056 4884 4064
rect 4892 4056 4900 4064
rect 4876 4016 4884 4024
rect 4814 4006 4822 4014
rect 4828 4006 4836 4014
rect 4842 4006 4850 4014
rect 5020 4256 5028 4264
rect 5052 4236 5060 4244
rect 5004 4196 5012 4204
rect 5084 4216 5092 4224
rect 5068 4196 5076 4204
rect 5116 4196 5124 4204
rect 5260 4636 5268 4644
rect 5500 5036 5508 5044
rect 5516 5036 5524 5044
rect 5548 5016 5556 5024
rect 5516 4996 5524 5004
rect 5532 4976 5540 4984
rect 5596 5016 5604 5024
rect 5836 5216 5844 5224
rect 5836 5176 5844 5184
rect 5756 5076 5764 5084
rect 5708 4976 5716 4984
rect 6252 5476 6260 5484
rect 6284 5376 6292 5384
rect 6380 5476 6388 5484
rect 6492 5476 6500 5484
rect 6380 5436 6388 5444
rect 6428 5436 6436 5444
rect 6350 5406 6358 5414
rect 6364 5406 6372 5414
rect 6378 5406 6386 5414
rect 6140 5336 6148 5344
rect 6220 5336 6228 5344
rect 6284 5336 6292 5344
rect 6316 5336 6324 5344
rect 5996 5316 6004 5324
rect 5948 5296 5956 5304
rect 6028 5256 6036 5264
rect 5948 5176 5956 5184
rect 6268 5316 6276 5324
rect 6172 5256 6180 5264
rect 6220 5296 6228 5304
rect 6268 5236 6276 5244
rect 6204 5196 6212 5204
rect 6204 5156 6212 5164
rect 6236 5156 6244 5164
rect 6236 5136 6244 5144
rect 6140 5116 6148 5124
rect 5916 5096 5924 5104
rect 5900 5056 5908 5064
rect 5788 5016 5796 5024
rect 5772 4996 5780 5004
rect 5404 4936 5412 4944
rect 5564 4936 5572 4944
rect 5644 4936 5652 4944
rect 5740 4936 5748 4944
rect 5356 4896 5364 4904
rect 5452 4916 5460 4924
rect 5676 4916 5684 4924
rect 5692 4916 5700 4924
rect 5756 4916 5764 4924
rect 5436 4896 5444 4904
rect 5452 4876 5460 4884
rect 5548 4876 5556 4884
rect 5468 4856 5476 4864
rect 5404 4836 5412 4844
rect 5340 4716 5348 4724
rect 5356 4716 5364 4724
rect 5388 4716 5396 4724
rect 5324 4696 5332 4704
rect 5324 4656 5332 4664
rect 5228 4556 5236 4564
rect 5388 4536 5396 4544
rect 5436 4756 5444 4764
rect 5452 4716 5460 4724
rect 5548 4856 5556 4864
rect 5580 4856 5588 4864
rect 5724 4896 5732 4904
rect 5756 4896 5764 4904
rect 5820 4856 5828 4864
rect 5708 4836 5716 4844
rect 5516 4756 5524 4764
rect 5532 4716 5540 4724
rect 5500 4696 5508 4704
rect 5516 4696 5524 4704
rect 5596 4696 5604 4704
rect 5628 4696 5636 4704
rect 5644 4676 5652 4684
rect 5676 4696 5684 4704
rect 5452 4656 5460 4664
rect 5484 4656 5492 4664
rect 5548 4656 5556 4664
rect 5500 4616 5508 4624
rect 5724 4676 5732 4684
rect 5740 4676 5748 4684
rect 5708 4656 5716 4664
rect 5692 4636 5700 4644
rect 5756 4636 5764 4644
rect 5500 4576 5508 4584
rect 5628 4576 5636 4584
rect 5660 4576 5668 4584
rect 5692 4576 5700 4584
rect 5548 4536 5556 4544
rect 5612 4536 5620 4544
rect 5404 4496 5412 4504
rect 5324 4476 5332 4484
rect 5292 4416 5300 4424
rect 5228 4396 5236 4404
rect 5820 4676 5828 4684
rect 5788 4656 5796 4664
rect 5788 4636 5796 4644
rect 5772 4616 5780 4624
rect 5772 4596 5780 4604
rect 5676 4556 5684 4564
rect 5756 4556 5764 4564
rect 5660 4536 5668 4544
rect 5724 4536 5732 4544
rect 5532 4516 5540 4524
rect 5564 4516 5572 4524
rect 5628 4516 5636 4524
rect 5580 4496 5588 4504
rect 5756 4516 5764 4524
rect 5724 4496 5732 4504
rect 5516 4476 5524 4484
rect 5564 4476 5572 4484
rect 5612 4476 5620 4484
rect 5420 4436 5428 4444
rect 5260 4296 5268 4304
rect 5308 4296 5316 4304
rect 5996 5016 6004 5024
rect 6028 4956 6036 4964
rect 5964 4936 5972 4944
rect 6060 4936 6068 4944
rect 6108 4936 6116 4944
rect 5932 4716 5940 4724
rect 5964 4716 5972 4724
rect 5852 4696 5860 4704
rect 5932 4696 5940 4704
rect 5948 4656 5956 4664
rect 5884 4616 5892 4624
rect 5868 4596 5876 4604
rect 5884 4556 5892 4564
rect 5884 4536 5892 4544
rect 5820 4516 5828 4524
rect 5884 4516 5892 4524
rect 5804 4416 5812 4424
rect 5932 4596 5940 4604
rect 6028 4776 6036 4784
rect 6044 4756 6052 4764
rect 6076 4736 6084 4744
rect 6012 4696 6020 4704
rect 5996 4596 6004 4604
rect 5948 4576 5956 4584
rect 6364 5376 6372 5384
rect 6316 5316 6324 5324
rect 6332 5316 6340 5324
rect 6332 5276 6340 5284
rect 6300 5236 6308 5244
rect 6348 5256 6356 5264
rect 6300 5156 6308 5164
rect 6332 5156 6340 5164
rect 6204 5096 6212 5104
rect 6220 5096 6228 5104
rect 6172 5076 6180 5084
rect 6460 5316 6468 5324
rect 6380 5296 6388 5304
rect 6364 5176 6372 5184
rect 6348 5136 6356 5144
rect 6300 5076 6308 5084
rect 6332 5076 6340 5084
rect 6412 5136 6420 5144
rect 6588 5376 6596 5384
rect 6524 5336 6532 5344
rect 6588 5336 6596 5344
rect 6524 5316 6532 5324
rect 6572 5316 6580 5324
rect 6476 5296 6484 5304
rect 6492 5296 6500 5304
rect 6444 5256 6452 5264
rect 6444 5196 6452 5204
rect 6460 5156 6468 5164
rect 6508 5156 6516 5164
rect 6540 5296 6548 5304
rect 6540 5256 6548 5264
rect 6652 5476 6660 5484
rect 6780 5496 6788 5504
rect 6716 5456 6724 5464
rect 6700 5436 6708 5444
rect 6748 5436 6756 5444
rect 6716 5396 6724 5404
rect 6796 5396 6804 5404
rect 6764 5376 6772 5384
rect 6732 5356 6740 5364
rect 6780 5356 6788 5364
rect 6796 5336 6804 5344
rect 6700 5316 6708 5324
rect 6620 5296 6628 5304
rect 6636 5276 6644 5284
rect 6940 5696 6948 5704
rect 7004 5696 7012 5704
rect 7020 5696 7028 5704
rect 6956 5676 6964 5684
rect 6972 5656 6980 5664
rect 6988 5636 6996 5644
rect 6876 5456 6884 5464
rect 7036 5436 7044 5444
rect 7004 5336 7012 5344
rect 7020 5336 7028 5344
rect 6988 5316 6996 5324
rect 6876 5296 6884 5304
rect 6828 5216 6836 5224
rect 6604 5156 6612 5164
rect 6572 5136 6580 5144
rect 6524 5116 6532 5124
rect 6428 5096 6436 5104
rect 6492 5096 6500 5104
rect 6476 5076 6484 5084
rect 6156 5036 6164 5044
rect 6380 5036 6388 5044
rect 6350 5006 6358 5014
rect 6364 5006 6372 5014
rect 6378 5006 6386 5014
rect 6284 4976 6292 4984
rect 6300 4936 6308 4944
rect 6220 4916 6228 4924
rect 6156 4856 6164 4864
rect 6220 4856 6228 4864
rect 6204 4836 6212 4844
rect 6204 4716 6212 4724
rect 6156 4696 6164 4704
rect 6156 4676 6164 4684
rect 6108 4636 6116 4644
rect 6140 4636 6148 4644
rect 6092 4556 6100 4564
rect 6316 4836 6324 4844
rect 6428 4916 6436 4924
rect 6428 4896 6436 4904
rect 6540 5076 6548 5084
rect 6492 4918 6500 4924
rect 6492 4916 6500 4918
rect 6460 4736 6468 4744
rect 6236 4716 6244 4724
rect 6316 4696 6324 4704
rect 6892 5102 6900 5104
rect 6892 5096 6900 5102
rect 6572 5036 6580 5044
rect 6636 5036 6644 5044
rect 7020 5296 7028 5304
rect 6732 5076 6740 5084
rect 6828 5076 6836 5084
rect 7100 5716 7108 5724
rect 7132 5716 7140 5724
rect 7148 5716 7156 5724
rect 7084 5696 7092 5704
rect 7196 5696 7204 5704
rect 7132 5676 7140 5684
rect 7148 5676 7156 5684
rect 7212 5676 7220 5684
rect 7100 5656 7108 5664
rect 7212 5656 7220 5664
rect 7132 5496 7140 5504
rect 7116 5476 7124 5484
rect 7084 5456 7092 5464
rect 7116 5456 7124 5464
rect 7068 5436 7076 5444
rect 7100 5396 7108 5404
rect 7132 5376 7140 5384
rect 7084 5336 7092 5344
rect 7068 5296 7076 5304
rect 7100 5296 7108 5304
rect 7068 5076 7076 5084
rect 7164 5516 7172 5524
rect 7324 5716 7332 5724
rect 7260 5696 7268 5704
rect 7276 5636 7284 5644
rect 7404 5576 7412 5584
rect 7276 5496 7284 5504
rect 7228 5476 7236 5484
rect 7260 5476 7268 5484
rect 7180 5456 7188 5464
rect 7244 5396 7252 5404
rect 7196 5356 7204 5364
rect 7276 5376 7284 5384
rect 7420 5536 7428 5544
rect 7340 5436 7348 5444
rect 7420 5436 7428 5444
rect 7148 5276 7156 5284
rect 7180 5316 7188 5324
rect 7164 5256 7172 5264
rect 7132 5156 7140 5164
rect 7164 5156 7172 5164
rect 7164 5136 7172 5144
rect 6956 5056 6964 5064
rect 6732 5036 6740 5044
rect 6764 5036 6772 5044
rect 6700 5016 6708 5024
rect 6572 4836 6580 4844
rect 6556 4716 6564 4724
rect 6620 4876 6628 4884
rect 6220 4676 6228 4684
rect 6284 4676 6292 4684
rect 6412 4676 6420 4684
rect 6396 4656 6404 4664
rect 6172 4636 6180 4644
rect 6364 4636 6372 4644
rect 6044 4536 6052 4544
rect 6350 4606 6358 4614
rect 6364 4606 6372 4614
rect 6378 4606 6386 4614
rect 6476 4656 6484 4664
rect 6508 4656 6516 4664
rect 6988 5016 6996 5024
rect 6764 4976 6772 4984
rect 6780 4936 6788 4944
rect 6668 4916 6676 4924
rect 6700 4916 6708 4924
rect 6652 4896 6660 4904
rect 6668 4876 6676 4884
rect 6796 4916 6804 4924
rect 6748 4876 6756 4884
rect 6684 4756 6692 4764
rect 6732 4756 6740 4764
rect 6652 4716 6660 4724
rect 6732 4716 6740 4724
rect 6860 4936 6868 4944
rect 6924 4936 6932 4944
rect 6828 4756 6836 4764
rect 6812 4716 6820 4724
rect 6700 4696 6708 4704
rect 6748 4696 6756 4704
rect 6796 4696 6804 4704
rect 6604 4676 6612 4684
rect 6636 4676 6644 4684
rect 6812 4676 6820 4684
rect 6924 4916 6932 4924
rect 6972 4916 6980 4924
rect 6876 4896 6884 4904
rect 6908 4896 6916 4904
rect 6956 4896 6964 4904
rect 6892 4876 6900 4884
rect 6924 4876 6932 4884
rect 6892 4756 6900 4764
rect 6844 4736 6852 4744
rect 6876 4736 6884 4744
rect 6908 4736 6916 4744
rect 7244 5336 7252 5344
rect 7292 5316 7300 5324
rect 7404 5376 7412 5384
rect 7356 5336 7364 5344
rect 7388 5316 7396 5324
rect 7404 5316 7412 5324
rect 7324 5296 7332 5304
rect 7468 5516 7476 5524
rect 7516 5476 7524 5484
rect 7452 5376 7460 5384
rect 7452 5316 7460 5324
rect 7228 5276 7236 5284
rect 7292 5276 7300 5284
rect 7436 5256 7444 5264
rect 7292 5156 7300 5164
rect 7388 5136 7396 5144
rect 7228 5076 7236 5084
rect 7196 5056 7204 5064
rect 7292 5076 7300 5084
rect 7052 5036 7060 5044
rect 7212 5036 7220 5044
rect 7244 5036 7252 5044
rect 7132 4976 7140 4984
rect 7036 4956 7044 4964
rect 7036 4936 7044 4944
rect 7260 4936 7268 4944
rect 6860 4716 6868 4724
rect 7116 4916 7124 4924
rect 7084 4876 7092 4884
rect 6956 4716 6964 4724
rect 6924 4696 6932 4704
rect 6956 4696 6964 4704
rect 7068 4756 7076 4764
rect 7036 4696 7044 4704
rect 7244 4918 7252 4924
rect 7244 4916 7252 4918
rect 7356 5056 7364 5064
rect 7404 5056 7412 5064
rect 7372 5036 7380 5044
rect 7324 5016 7332 5024
rect 7404 5016 7412 5024
rect 7388 4996 7396 5004
rect 7276 4776 7284 4784
rect 7292 4716 7300 4724
rect 7404 4696 7412 4704
rect 7436 4716 7444 4724
rect 7084 4676 7092 4684
rect 7132 4676 7140 4684
rect 7180 4676 7188 4684
rect 6540 4656 6548 4664
rect 6572 4656 6580 4664
rect 6796 4656 6804 4664
rect 6988 4656 6996 4664
rect 7100 4656 7108 4664
rect 7148 4656 7156 4664
rect 6524 4636 6532 4644
rect 6620 4636 6628 4644
rect 6444 4576 6452 4584
rect 6620 4576 6628 4584
rect 6796 4576 6804 4584
rect 6284 4556 6292 4564
rect 6492 4556 6500 4564
rect 6524 4556 6532 4564
rect 6636 4556 6644 4564
rect 6700 4556 6708 4564
rect 6252 4536 6260 4544
rect 6604 4536 6612 4544
rect 5836 4396 5844 4404
rect 5580 4356 5588 4364
rect 5756 4356 5764 4364
rect 5884 4356 5892 4364
rect 5468 4336 5476 4344
rect 5708 4336 5716 4344
rect 5740 4336 5748 4344
rect 5868 4336 5876 4344
rect 5612 4296 5620 4304
rect 5660 4296 5668 4304
rect 5724 4296 5732 4304
rect 5212 4256 5220 4264
rect 5244 4256 5252 4264
rect 5196 4236 5204 4244
rect 5244 4216 5252 4224
rect 5324 4196 5332 4204
rect 5180 4176 5188 4184
rect 5228 4176 5236 4184
rect 5340 4156 5348 4164
rect 5036 4116 5044 4124
rect 5116 4116 5124 4124
rect 5020 4096 5028 4104
rect 5100 4096 5108 4104
rect 5196 4096 5204 4104
rect 5036 4076 5044 4084
rect 5068 4076 5076 4084
rect 5084 4076 5092 4084
rect 4956 3936 4964 3944
rect 4988 3936 4996 3944
rect 4796 3856 4804 3864
rect 4780 3796 4788 3804
rect 4748 3756 4756 3764
rect 4780 3716 4788 3724
rect 4556 3696 4564 3704
rect 4604 3676 4612 3684
rect 4604 3636 4612 3644
rect 4636 3696 4644 3704
rect 4668 3696 4676 3704
rect 4764 3696 4772 3704
rect 4828 3716 4836 3724
rect 4876 3856 4884 3864
rect 4924 3836 4932 3844
rect 4940 3836 4948 3844
rect 4956 3836 4964 3844
rect 4876 3816 4884 3824
rect 4860 3656 4868 3664
rect 4812 3636 4820 3644
rect 4524 3576 4532 3584
rect 4620 3576 4628 3584
rect 4814 3606 4822 3614
rect 4828 3606 4836 3614
rect 4842 3606 4850 3614
rect 4748 3596 4756 3604
rect 4444 3556 4452 3564
rect 4684 3556 4692 3564
rect 4508 3536 4516 3544
rect 4524 3536 4532 3544
rect 4364 3496 4372 3504
rect 4396 3496 4404 3504
rect 4444 3496 4452 3504
rect 4364 3476 4372 3484
rect 4556 3516 4564 3524
rect 4620 3516 4628 3524
rect 4828 3516 4836 3524
rect 4588 3496 4596 3504
rect 4700 3496 4708 3504
rect 4492 3476 4500 3484
rect 4428 3436 4436 3444
rect 4476 3356 4484 3364
rect 4300 3336 4308 3344
rect 4348 3340 4356 3344
rect 4348 3336 4356 3340
rect 4284 3316 4292 3324
rect 3916 3296 3924 3304
rect 3980 3296 3988 3304
rect 4060 3296 4068 3304
rect 4188 3296 4196 3304
rect 4252 3296 4260 3304
rect 3708 3276 3716 3284
rect 3836 3276 3844 3284
rect 3788 3156 3796 3164
rect 3580 3136 3588 3144
rect 3612 3136 3620 3144
rect 3644 3136 3652 3144
rect 3692 3136 3700 3144
rect 3564 3116 3572 3124
rect 3420 3076 3428 3084
rect 3452 3076 3460 3084
rect 3340 3056 3348 3064
rect 3180 2976 3188 2984
rect 3148 2956 3156 2964
rect 2924 2776 2932 2784
rect 2956 2776 2964 2784
rect 2476 2696 2484 2704
rect 2620 2676 2628 2684
rect 2492 2636 2500 2644
rect 2556 2636 2564 2644
rect 2636 2636 2644 2644
rect 2524 2616 2532 2624
rect 2796 2696 2804 2704
rect 2988 2696 2996 2704
rect 2700 2676 2708 2684
rect 2732 2656 2740 2664
rect 2668 2616 2676 2624
rect 2860 2596 2868 2604
rect 2588 2556 2596 2564
rect 3052 2918 3060 2924
rect 3052 2916 3060 2918
rect 3196 2836 3204 2844
rect 3278 3006 3286 3014
rect 3292 3006 3300 3014
rect 3306 3006 3314 3014
rect 3516 3056 3524 3064
rect 3468 2996 3476 3004
rect 3372 2976 3380 2984
rect 3356 2956 3364 2964
rect 3404 2956 3412 2964
rect 3324 2936 3332 2944
rect 3452 2916 3460 2924
rect 3740 3116 3748 3124
rect 4204 3256 4212 3264
rect 4204 3196 4212 3204
rect 3884 3136 3892 3144
rect 3852 3116 3860 3124
rect 3548 3056 3556 3064
rect 3548 3016 3556 3024
rect 3532 2996 3540 3004
rect 3484 2976 3492 2984
rect 3500 2976 3508 2984
rect 3532 2976 3540 2984
rect 3628 3076 3636 3084
rect 3788 3076 3796 3084
rect 3836 3076 3844 3084
rect 3724 3056 3732 3064
rect 3980 3116 3988 3124
rect 4252 3176 4260 3184
rect 4044 3076 4052 3084
rect 4076 3076 4084 3084
rect 4236 3076 4244 3084
rect 3804 3056 3812 3064
rect 3852 3056 3860 3064
rect 3884 3056 3892 3064
rect 3772 3016 3780 3024
rect 3644 2976 3652 2984
rect 3676 2976 3684 2984
rect 3756 2976 3764 2984
rect 3484 2936 3492 2944
rect 3516 2936 3524 2944
rect 3324 2876 3332 2884
rect 3660 2956 3668 2964
rect 3772 2956 3780 2964
rect 3420 2856 3428 2864
rect 3548 2876 3556 2884
rect 3804 2936 3812 2944
rect 3628 2916 3636 2924
rect 3884 3016 3892 3024
rect 3900 2996 3908 3004
rect 4044 2996 4052 3004
rect 3980 2956 3988 2964
rect 3820 2916 3828 2924
rect 3852 2916 3860 2924
rect 3868 2916 3876 2924
rect 3596 2896 3604 2904
rect 3820 2896 3828 2904
rect 3580 2856 3588 2864
rect 3516 2836 3524 2844
rect 3116 2776 3124 2784
rect 3052 2702 3060 2704
rect 3052 2696 3060 2702
rect 3244 2736 3252 2744
rect 3196 2716 3204 2724
rect 3180 2696 3188 2704
rect 3388 2702 3396 2704
rect 3388 2696 3396 2702
rect 3452 2696 3460 2704
rect 3484 2696 3492 2704
rect 3164 2656 3172 2664
rect 3196 2656 3204 2664
rect 3244 2656 3252 2664
rect 2956 2636 2964 2644
rect 2972 2596 2980 2604
rect 3100 2596 3108 2604
rect 2908 2576 2916 2584
rect 2876 2556 2884 2564
rect 3084 2576 3092 2584
rect 3278 2606 3286 2614
rect 3292 2606 3300 2614
rect 3306 2606 3314 2614
rect 3244 2576 3252 2584
rect 3116 2556 3124 2564
rect 3228 2556 3236 2564
rect 2476 2536 2484 2544
rect 2572 2536 2580 2544
rect 2428 2496 2436 2504
rect 2460 2376 2468 2384
rect 2492 2516 2500 2524
rect 2540 2516 2548 2524
rect 2684 2496 2692 2504
rect 2636 2356 2644 2364
rect 2908 2516 2916 2524
rect 2892 2496 2900 2504
rect 2988 2496 2996 2504
rect 2956 2476 2964 2484
rect 2796 2456 2804 2464
rect 2876 2376 2884 2384
rect 2924 2356 2932 2364
rect 2844 2336 2852 2344
rect 2892 2336 2900 2344
rect 3036 2516 3044 2524
rect 3132 2516 3140 2524
rect 3212 2536 3220 2544
rect 3164 2516 3172 2524
rect 3260 2556 3268 2564
rect 3308 2536 3316 2544
rect 3356 2536 3364 2544
rect 3180 2496 3188 2504
rect 3196 2476 3204 2484
rect 3276 2476 3284 2484
rect 3356 2476 3364 2484
rect 3052 2456 3060 2464
rect 3180 2396 3188 2404
rect 3020 2336 3028 2344
rect 2732 2316 2740 2324
rect 2796 2316 2804 2324
rect 2988 2316 2996 2324
rect 3148 2316 3156 2324
rect 2620 2296 2628 2304
rect 2668 2296 2676 2304
rect 2476 2276 2484 2284
rect 2380 2256 2388 2264
rect 2572 2256 2580 2264
rect 2636 2256 2644 2264
rect 2588 2236 2596 2244
rect 2636 2236 2644 2244
rect 2364 2216 2372 2224
rect 2572 2216 2580 2224
rect 2428 2176 2436 2184
rect 2380 2136 2388 2144
rect 2332 1956 2340 1964
rect 2316 1936 2324 1944
rect 2556 2136 2564 2144
rect 2620 2196 2628 2204
rect 2652 2216 2660 2224
rect 2700 2256 2708 2264
rect 2652 2196 2660 2204
rect 2684 2196 2692 2204
rect 2588 2116 2596 2124
rect 2572 2076 2580 2084
rect 2684 2176 2692 2184
rect 2796 2296 2804 2304
rect 2844 2296 2852 2304
rect 2748 2276 2756 2284
rect 2860 2276 2868 2284
rect 2812 2236 2820 2244
rect 2796 2216 2804 2224
rect 2732 2156 2740 2164
rect 2764 2156 2772 2164
rect 2684 2096 2692 2104
rect 2860 2196 2868 2204
rect 3004 2296 3012 2304
rect 2956 2256 2964 2264
rect 3036 2276 3044 2284
rect 3100 2276 3108 2284
rect 3148 2276 3156 2284
rect 2844 2176 2852 2184
rect 3052 2256 3060 2264
rect 3164 2256 3172 2264
rect 3276 2336 3284 2344
rect 3340 2296 3348 2304
rect 3388 2656 3396 2664
rect 3420 2656 3428 2664
rect 3452 2636 3460 2644
rect 3452 2616 3460 2624
rect 3436 2556 3444 2564
rect 3500 2536 3508 2544
rect 3468 2516 3476 2524
rect 3420 2496 3428 2504
rect 3484 2496 3492 2504
rect 3468 2476 3476 2484
rect 3404 2302 3412 2304
rect 3404 2296 3412 2302
rect 3468 2296 3476 2304
rect 3278 2206 3286 2214
rect 3292 2206 3300 2214
rect 3306 2206 3314 2214
rect 2988 2156 2996 2164
rect 3036 2156 3044 2164
rect 3068 2156 3076 2164
rect 3164 2176 3172 2184
rect 3500 2236 3508 2244
rect 3996 2936 4004 2944
rect 3916 2896 3924 2904
rect 4172 2976 4180 2984
rect 4092 2936 4100 2944
rect 4284 2956 4292 2964
rect 3948 2896 3956 2904
rect 3996 2896 4004 2904
rect 4076 2856 4084 2864
rect 3932 2836 3940 2844
rect 3548 2736 3556 2744
rect 3788 2736 3796 2744
rect 3884 2736 3892 2744
rect 3724 2716 3732 2724
rect 3580 2696 3588 2704
rect 3692 2676 3700 2684
rect 3596 2656 3604 2664
rect 3692 2656 3700 2664
rect 3532 2576 3540 2584
rect 3596 2536 3604 2544
rect 3532 2476 3540 2484
rect 3580 2476 3588 2484
rect 3660 2476 3668 2484
rect 4140 2916 4148 2924
rect 4060 2736 4068 2744
rect 3836 2676 3844 2684
rect 3756 2656 3764 2664
rect 3836 2656 3844 2664
rect 3724 2616 3732 2624
rect 3708 2576 3716 2584
rect 3788 2576 3796 2584
rect 3804 2536 3812 2544
rect 3820 2536 3828 2544
rect 3708 2516 3716 2524
rect 3548 2296 3556 2304
rect 3708 2296 3716 2304
rect 3756 2296 3764 2304
rect 3804 2296 3812 2304
rect 3724 2276 3732 2284
rect 3532 2216 3540 2224
rect 3692 2156 3700 2164
rect 2748 2136 2756 2144
rect 2764 2136 2772 2144
rect 2924 2136 2932 2144
rect 2972 2136 2980 2144
rect 3676 2136 3684 2144
rect 2892 2116 2900 2124
rect 3020 2116 3028 2124
rect 3308 2118 3316 2124
rect 3308 2116 3316 2118
rect 3468 2116 3476 2124
rect 2764 2096 2772 2104
rect 2812 2096 2820 2104
rect 3164 2096 3172 2104
rect 3420 2096 3428 2104
rect 2716 2076 2724 2084
rect 2780 2076 2788 2084
rect 2860 2076 2868 2084
rect 2940 2076 2948 2084
rect 3148 2076 3156 2084
rect 2812 2056 2820 2064
rect 2700 1996 2708 2004
rect 2764 1996 2772 2004
rect 2492 1956 2500 1964
rect 2556 1956 2564 1964
rect 2444 1936 2452 1944
rect 2396 1916 2404 1924
rect 2332 1876 2340 1884
rect 2396 1896 2404 1904
rect 2524 1896 2532 1904
rect 2380 1876 2388 1884
rect 2524 1876 2532 1884
rect 2572 1876 2580 1884
rect 2668 1876 2676 1884
rect 2684 1876 2692 1884
rect 2748 1876 2756 1884
rect 2588 1856 2596 1864
rect 2652 1856 2660 1864
rect 2540 1796 2548 1804
rect 2428 1776 2436 1784
rect 2492 1776 2500 1784
rect 2508 1776 2516 1784
rect 2396 1756 2404 1764
rect 2604 1816 2612 1824
rect 2588 1776 2596 1784
rect 2332 1696 2340 1704
rect 2348 1636 2356 1644
rect 2284 1516 2292 1524
rect 2172 1496 2180 1504
rect 2172 1396 2180 1404
rect 2284 1496 2292 1504
rect 2316 1496 2324 1504
rect 2444 1676 2452 1684
rect 2700 1856 2708 1864
rect 2716 1756 2724 1764
rect 2636 1736 2644 1744
rect 2652 1736 2660 1744
rect 2604 1676 2612 1684
rect 2668 1676 2676 1684
rect 2700 1736 2708 1744
rect 2796 1956 2804 1964
rect 2828 1976 2836 1984
rect 2876 1976 2884 1984
rect 2812 1876 2820 1884
rect 3100 1936 3108 1944
rect 3356 2076 3364 2084
rect 3068 1916 3076 1924
rect 3132 1916 3140 1924
rect 2972 1896 2980 1904
rect 3036 1896 3044 1904
rect 2908 1876 2916 1884
rect 2812 1856 2820 1864
rect 3004 1856 3012 1864
rect 2780 1836 2788 1844
rect 2780 1816 2788 1824
rect 2716 1696 2724 1704
rect 2732 1696 2740 1704
rect 2540 1656 2548 1664
rect 2684 1656 2692 1664
rect 2460 1636 2468 1644
rect 2684 1636 2692 1644
rect 2588 1576 2596 1584
rect 2668 1516 2676 1524
rect 2300 1476 2308 1484
rect 2556 1476 2564 1484
rect 2268 1436 2276 1444
rect 2252 1416 2260 1424
rect 2300 1416 2308 1424
rect 2492 1376 2500 1384
rect 2124 1336 2132 1344
rect 2076 1316 2084 1324
rect 2044 1196 2052 1204
rect 2044 1176 2052 1184
rect 2028 1156 2036 1164
rect 2012 1056 2020 1064
rect 2044 1056 2052 1064
rect 2012 1036 2020 1044
rect 2012 976 2020 984
rect 1932 936 1940 944
rect 1980 896 1988 904
rect 2092 1096 2100 1104
rect 2220 1356 2228 1364
rect 2252 1356 2260 1364
rect 2332 1356 2340 1364
rect 2188 1336 2196 1344
rect 2156 1296 2164 1304
rect 2236 1276 2244 1284
rect 2220 1216 2228 1224
rect 2140 1196 2148 1204
rect 2124 1136 2132 1144
rect 2156 1096 2164 1104
rect 2204 1096 2212 1104
rect 2332 1316 2340 1324
rect 2348 1236 2356 1244
rect 2316 1156 2324 1164
rect 2332 1136 2340 1144
rect 2316 1116 2324 1124
rect 2412 1316 2420 1324
rect 2396 1196 2404 1204
rect 2412 1176 2420 1184
rect 2396 1156 2404 1164
rect 2364 1136 2372 1144
rect 2492 1316 2500 1324
rect 2748 1616 2756 1624
rect 2908 1836 2916 1844
rect 2828 1796 2836 1804
rect 2844 1756 2852 1764
rect 2812 1716 2820 1724
rect 2780 1636 2788 1644
rect 2892 1816 2900 1824
rect 2876 1776 2884 1784
rect 2892 1676 2900 1684
rect 2860 1596 2868 1604
rect 2764 1576 2772 1584
rect 2940 1796 2948 1804
rect 2924 1736 2932 1744
rect 2956 1676 2964 1684
rect 2988 1636 2996 1644
rect 3276 2016 3284 2024
rect 3228 1936 3236 1944
rect 3260 1916 3268 1924
rect 3084 1896 3092 1904
rect 3180 1896 3188 1904
rect 3132 1876 3140 1884
rect 3196 1876 3204 1884
rect 3180 1856 3188 1864
rect 3500 2096 3508 2104
rect 3452 2016 3460 2024
rect 3356 1956 3364 1964
rect 3340 1916 3348 1924
rect 3260 1876 3268 1884
rect 3052 1836 3060 1844
rect 3212 1836 3220 1844
rect 3244 1816 3252 1824
rect 3278 1806 3286 1814
rect 3292 1806 3300 1814
rect 3306 1806 3314 1814
rect 3068 1776 3076 1784
rect 3244 1776 3252 1784
rect 3324 1776 3332 1784
rect 3036 1756 3044 1764
rect 3052 1756 3060 1764
rect 3196 1756 3204 1764
rect 3276 1756 3284 1764
rect 3388 1856 3396 1864
rect 3372 1836 3380 1844
rect 3356 1756 3364 1764
rect 3372 1756 3380 1764
rect 3468 1956 3476 1964
rect 3436 1876 3444 1884
rect 3452 1796 3460 1804
rect 3436 1776 3444 1784
rect 3148 1736 3156 1744
rect 3180 1736 3188 1744
rect 3212 1736 3220 1744
rect 3260 1736 3268 1744
rect 3356 1736 3364 1744
rect 3404 1736 3412 1744
rect 3420 1736 3428 1744
rect 3100 1716 3108 1724
rect 3020 1676 3028 1684
rect 3020 1656 3028 1664
rect 3148 1696 3156 1704
rect 3164 1696 3172 1704
rect 3212 1696 3220 1704
rect 3260 1696 3268 1704
rect 3404 1656 3412 1664
rect 3116 1636 3124 1644
rect 3212 1636 3220 1644
rect 3452 1636 3460 1644
rect 3132 1616 3140 1624
rect 3260 1536 3268 1544
rect 3004 1516 3012 1524
rect 3228 1516 3236 1524
rect 2828 1496 2836 1504
rect 3100 1496 3108 1504
rect 3356 1496 3364 1504
rect 3468 1496 3476 1504
rect 2716 1476 2724 1484
rect 2860 1476 2868 1484
rect 3052 1476 3060 1484
rect 3244 1476 3252 1484
rect 3420 1476 3428 1484
rect 2460 1176 2468 1184
rect 2476 1156 2484 1164
rect 2412 1116 2420 1124
rect 2428 1116 2436 1124
rect 2364 1096 2372 1104
rect 2620 1276 2628 1284
rect 2668 1276 2676 1284
rect 2572 1236 2580 1244
rect 2636 1236 2644 1244
rect 2508 1136 2516 1144
rect 2588 1216 2596 1224
rect 2412 1096 2420 1104
rect 2492 1096 2500 1104
rect 2540 1096 2548 1104
rect 2108 1076 2116 1084
rect 2140 1076 2148 1084
rect 2204 1076 2212 1084
rect 2332 1076 2340 1084
rect 2396 1076 2404 1084
rect 2188 1056 2196 1064
rect 2060 1036 2068 1044
rect 2380 1056 2388 1064
rect 2492 1056 2500 1064
rect 2252 1036 2260 1044
rect 2300 1036 2308 1044
rect 2444 1036 2452 1044
rect 2220 996 2228 1004
rect 2204 976 2212 984
rect 2524 1016 2532 1024
rect 2428 936 2436 944
rect 2140 918 2148 924
rect 2140 916 2148 918
rect 2172 916 2180 924
rect 2124 896 2132 904
rect 2172 896 2180 904
rect 2060 816 2068 824
rect 1916 702 1924 704
rect 1916 696 1924 702
rect 2348 756 2356 764
rect 2204 736 2212 744
rect 2268 736 2276 744
rect 1852 656 1860 664
rect 1836 636 1844 644
rect 1596 616 1604 624
rect 1676 616 1684 624
rect 1980 656 1988 664
rect 2220 716 2228 724
rect 2284 716 2292 724
rect 2332 716 2340 724
rect 2236 676 2244 684
rect 1580 576 1588 584
rect 1388 556 1396 564
rect 1228 456 1236 464
rect 2060 596 2068 604
rect 2492 756 2500 764
rect 2380 716 2388 724
rect 2412 716 2420 724
rect 2476 716 2484 724
rect 2268 676 2276 684
rect 2332 676 2340 684
rect 2188 576 2196 584
rect 1564 556 1572 564
rect 1644 556 1652 564
rect 2060 556 2068 564
rect 2124 556 2132 564
rect 2236 556 2244 564
rect 1532 536 1540 544
rect 1580 536 1588 544
rect 1868 536 1876 544
rect 1836 516 1844 524
rect 1564 496 1572 504
rect 1644 496 1652 504
rect 1676 496 1684 504
rect 1644 476 1652 484
rect 1692 476 1700 484
rect 1308 316 1316 324
rect 1742 406 1750 414
rect 1756 406 1764 414
rect 1770 406 1778 414
rect 1420 336 1428 344
rect 1564 336 1572 344
rect 1580 336 1588 344
rect 1740 336 1748 344
rect 1452 316 1460 324
rect 1548 316 1556 324
rect 1676 316 1684 324
rect 1708 316 1716 324
rect 1756 316 1764 324
rect 1148 276 1156 284
rect 1244 276 1252 284
rect 1340 276 1348 284
rect 940 256 948 264
rect 892 196 900 204
rect 892 136 900 144
rect 940 136 948 144
rect 1068 256 1076 264
rect 1164 256 1172 264
rect 1196 256 1204 264
rect 1308 216 1316 224
rect 1196 156 1204 164
rect 1388 216 1396 224
rect 1052 136 1060 144
rect 956 116 964 124
rect 1148 116 1156 124
rect 1260 116 1268 124
rect 1324 118 1332 124
rect 1324 116 1332 118
rect 1420 116 1428 124
rect 412 96 420 104
rect 748 96 756 104
rect 876 96 884 104
rect 1148 96 1156 104
rect 1676 296 1684 304
rect 1500 256 1508 264
rect 1532 236 1540 244
rect 1628 256 1636 264
rect 1612 236 1620 244
rect 1692 276 1700 284
rect 1692 256 1700 264
rect 1724 256 1732 264
rect 1628 216 1636 224
rect 1516 156 1524 164
rect 1532 156 1540 164
rect 1644 156 1652 164
rect 1676 156 1684 164
rect 1612 136 1620 144
rect 1580 116 1588 124
rect 1708 156 1716 164
rect 1996 536 2004 544
rect 2108 536 2116 544
rect 2316 656 2324 664
rect 2284 636 2292 644
rect 2284 616 2292 624
rect 2268 536 2276 544
rect 2428 696 2436 704
rect 2444 696 2452 704
rect 2476 696 2484 704
rect 2604 1176 2612 1184
rect 2620 1136 2628 1144
rect 2684 1136 2692 1144
rect 2652 1096 2660 1104
rect 3356 1436 3364 1444
rect 3278 1406 3286 1414
rect 3292 1406 3300 1414
rect 3306 1406 3314 1414
rect 3388 1376 3396 1384
rect 2876 1356 2884 1364
rect 2908 1356 2916 1364
rect 2892 1336 2900 1344
rect 3100 1336 3108 1344
rect 3036 1318 3044 1324
rect 3036 1316 3044 1318
rect 3132 1316 3140 1324
rect 3068 1296 3076 1304
rect 3228 1316 3236 1324
rect 3356 1316 3364 1324
rect 3452 1336 3460 1344
rect 3212 1296 3220 1304
rect 3388 1296 3396 1304
rect 3404 1296 3412 1304
rect 3436 1296 3444 1304
rect 3596 2116 3604 2124
rect 3660 2116 3668 2124
rect 3628 2096 3636 2104
rect 3532 2076 3540 2084
rect 3660 2016 3668 2024
rect 3644 1996 3652 2004
rect 3820 2256 3828 2264
rect 3868 2540 3876 2544
rect 3868 2536 3876 2540
rect 3884 2536 3892 2544
rect 4012 2616 4020 2624
rect 3964 2556 3972 2564
rect 3932 2536 3940 2544
rect 3900 2516 3908 2524
rect 4124 2856 4132 2864
rect 4124 2836 4132 2844
rect 4172 2676 4180 2684
rect 4236 2936 4244 2944
rect 4364 3316 4372 3324
rect 4460 3316 4468 3324
rect 4332 3056 4340 3064
rect 4316 2936 4324 2944
rect 4364 2856 4372 2864
rect 4300 2816 4308 2824
rect 4364 2796 4372 2804
rect 4204 2776 4212 2784
rect 4236 2756 4244 2764
rect 4268 2716 4276 2724
rect 4092 2596 4100 2604
rect 4108 2596 4116 2604
rect 4028 2576 4036 2584
rect 4076 2576 4084 2584
rect 4140 2576 4148 2584
rect 4220 2676 4228 2684
rect 4284 2676 4292 2684
rect 4556 3476 4564 3484
rect 4524 3236 4532 3244
rect 4636 3476 4644 3484
rect 4796 3496 4804 3504
rect 4812 3476 4820 3484
rect 4748 3456 4756 3464
rect 4796 3436 4804 3444
rect 4668 3416 4676 3424
rect 4684 3396 4692 3404
rect 4748 3396 4756 3404
rect 4620 3376 4628 3384
rect 4716 3356 4724 3364
rect 4828 3416 4836 3424
rect 4620 3336 4628 3344
rect 4812 3336 4820 3344
rect 4604 3316 4612 3324
rect 4732 3316 4740 3324
rect 4780 3316 4788 3324
rect 4732 3276 4740 3284
rect 4780 3236 4788 3244
rect 4814 3206 4822 3214
rect 4828 3206 4836 3214
rect 4842 3206 4850 3214
rect 4972 3816 4980 3824
rect 4972 3776 4980 3784
rect 5052 3816 5060 3824
rect 4988 3736 4996 3744
rect 5068 3736 5076 3744
rect 4924 3716 4932 3724
rect 4892 3696 4900 3704
rect 4908 3656 4916 3664
rect 4940 3576 4948 3584
rect 4956 3516 4964 3524
rect 4892 3496 4900 3504
rect 4908 3436 4916 3444
rect 4956 3436 4964 3444
rect 4972 3436 4980 3444
rect 4956 3376 4964 3384
rect 4940 3356 4948 3364
rect 4892 3336 4900 3344
rect 4972 3296 4980 3304
rect 5020 3656 5028 3664
rect 5164 3936 5172 3944
rect 5132 3876 5140 3884
rect 5292 4116 5300 4124
rect 5212 4016 5220 4024
rect 5228 4016 5236 4024
rect 5356 4136 5364 4144
rect 5372 4136 5380 4144
rect 5452 4196 5460 4204
rect 5468 4176 5476 4184
rect 5356 4116 5364 4124
rect 5388 4116 5396 4124
rect 5420 4116 5428 4124
rect 5308 4096 5316 4104
rect 5228 3996 5236 4004
rect 5276 3996 5284 4004
rect 5260 3936 5268 3944
rect 5372 4056 5380 4064
rect 5452 3956 5460 3964
rect 5340 3936 5348 3944
rect 5372 3936 5380 3944
rect 5484 3936 5492 3944
rect 5452 3916 5460 3924
rect 5180 3896 5188 3904
rect 5196 3896 5204 3904
rect 5228 3896 5236 3904
rect 5260 3896 5268 3904
rect 5404 3896 5412 3904
rect 5100 3756 5108 3764
rect 5292 3876 5300 3884
rect 5308 3876 5316 3884
rect 5292 3856 5300 3864
rect 5548 4276 5556 4284
rect 5708 4276 5716 4284
rect 5596 4236 5604 4244
rect 5644 4236 5652 4244
rect 5596 4216 5604 4224
rect 5516 4156 5524 4164
rect 5692 4156 5700 4164
rect 5644 4136 5652 4144
rect 5612 4116 5620 4124
rect 5788 4296 5796 4304
rect 5756 4276 5764 4284
rect 5804 4276 5812 4284
rect 5788 4256 5796 4264
rect 5868 4276 5876 4284
rect 5964 4336 5972 4344
rect 6028 4336 6036 4344
rect 5980 4276 5988 4284
rect 5900 4256 5908 4264
rect 5996 4256 6004 4264
rect 5836 4236 5844 4244
rect 5820 4216 5828 4224
rect 5868 4216 5876 4224
rect 5932 4216 5940 4224
rect 5852 4196 5860 4204
rect 5756 4176 5764 4184
rect 5852 4176 5860 4184
rect 5740 4156 5748 4164
rect 5756 4156 5764 4164
rect 5820 4156 5828 4164
rect 6012 4156 6020 4164
rect 5868 4136 5876 4144
rect 6220 4516 6228 4524
rect 6540 4516 6548 4524
rect 6204 4496 6212 4504
rect 6284 4496 6292 4504
rect 6412 4496 6420 4504
rect 6060 4476 6068 4484
rect 6108 4476 6116 4484
rect 6124 4456 6132 4464
rect 6556 4496 6564 4504
rect 6524 4476 6532 4484
rect 6684 4516 6692 4524
rect 6652 4496 6660 4504
rect 6764 4536 6772 4544
rect 6780 4536 6788 4544
rect 6828 4556 6836 4564
rect 6828 4536 6836 4544
rect 6908 4536 6916 4544
rect 6668 4476 6676 4484
rect 6748 4476 6756 4484
rect 6748 4436 6756 4444
rect 6300 4356 6308 4364
rect 6076 4336 6084 4344
rect 6124 4336 6132 4344
rect 6156 4336 6164 4344
rect 6204 4316 6212 4324
rect 6236 4316 6244 4324
rect 6284 4316 6292 4324
rect 6076 4296 6084 4304
rect 6076 4176 6084 4184
rect 6172 4276 6180 4284
rect 6140 4256 6148 4264
rect 6140 4216 6148 4224
rect 6204 4256 6212 4264
rect 6188 4236 6196 4244
rect 6316 4316 6324 4324
rect 6348 4316 6356 4324
rect 6524 4316 6532 4324
rect 6380 4296 6388 4304
rect 6444 4276 6452 4284
rect 6316 4256 6324 4264
rect 6412 4256 6420 4264
rect 6684 4336 6692 4344
rect 6748 4336 6756 4344
rect 6796 4336 6804 4344
rect 6604 4296 6612 4304
rect 6700 4296 6708 4304
rect 6716 4276 6724 4284
rect 6428 4236 6436 4244
rect 6252 4216 6260 4224
rect 6204 4196 6212 4204
rect 6188 4176 6196 4184
rect 6044 4136 6052 4144
rect 5772 4116 5780 4124
rect 6076 4116 6084 4124
rect 5564 4096 5572 4104
rect 5660 4096 5668 4104
rect 5692 4096 5700 4104
rect 5724 4096 5732 4104
rect 5628 4016 5636 4024
rect 5612 3996 5620 4004
rect 5516 3916 5524 3924
rect 5452 3876 5460 3884
rect 5388 3776 5396 3784
rect 5260 3756 5268 3764
rect 5308 3756 5316 3764
rect 5324 3756 5332 3764
rect 5196 3716 5204 3724
rect 5420 3856 5428 3864
rect 5820 4056 5828 4064
rect 5820 4016 5828 4024
rect 5660 3996 5668 4004
rect 5884 3996 5892 4004
rect 5852 3936 5860 3944
rect 5868 3936 5876 3944
rect 5948 3936 5956 3944
rect 5708 3916 5716 3924
rect 5740 3916 5748 3924
rect 5804 3916 5812 3924
rect 5836 3916 5844 3924
rect 5644 3896 5652 3904
rect 5692 3896 5700 3904
rect 5740 3896 5748 3904
rect 5756 3896 5764 3904
rect 5788 3876 5796 3884
rect 5932 3896 5940 3904
rect 5996 3896 6004 3904
rect 6028 3896 6036 3904
rect 6060 3902 6068 3904
rect 6060 3896 6068 3902
rect 5900 3876 5908 3884
rect 5980 3876 5988 3884
rect 5628 3856 5636 3864
rect 5756 3856 5764 3864
rect 5852 3856 5860 3864
rect 5900 3856 5908 3864
rect 5884 3836 5892 3844
rect 5788 3816 5796 3824
rect 5868 3796 5876 3804
rect 5420 3756 5428 3764
rect 5452 3756 5460 3764
rect 5292 3656 5300 3664
rect 5180 3576 5188 3584
rect 5612 3716 5620 3724
rect 5436 3616 5444 3624
rect 5436 3596 5444 3604
rect 5500 3596 5508 3604
rect 5292 3556 5300 3564
rect 5340 3556 5348 3564
rect 5372 3536 5380 3544
rect 5004 3516 5012 3524
rect 5260 3516 5268 3524
rect 5036 3496 5044 3504
rect 5196 3496 5204 3504
rect 5228 3496 5236 3504
rect 5100 3476 5108 3484
rect 5036 3456 5044 3464
rect 5084 3456 5092 3464
rect 5052 3436 5060 3444
rect 5004 3356 5012 3364
rect 5020 3356 5028 3364
rect 5052 3276 5060 3284
rect 4988 3256 4996 3264
rect 5292 3496 5300 3504
rect 5276 3476 5284 3484
rect 5404 3516 5412 3524
rect 5420 3516 5428 3524
rect 5500 3516 5508 3524
rect 5516 3516 5524 3524
rect 5340 3496 5348 3504
rect 5212 3456 5220 3464
rect 5324 3456 5332 3464
rect 5340 3456 5348 3464
rect 5196 3416 5204 3424
rect 5404 3496 5412 3504
rect 5452 3496 5460 3504
rect 5484 3496 5492 3504
rect 5516 3496 5524 3504
rect 5372 3476 5380 3484
rect 5420 3456 5428 3464
rect 5356 3416 5364 3424
rect 5260 3396 5268 3404
rect 5324 3396 5332 3404
rect 5100 3376 5108 3384
rect 5180 3376 5188 3384
rect 5084 3336 5092 3344
rect 5148 3336 5156 3344
rect 5164 3336 5172 3344
rect 5132 3316 5140 3324
rect 5356 3376 5364 3384
rect 5324 3356 5332 3364
rect 5228 3336 5236 3344
rect 5164 3296 5172 3304
rect 5052 3236 5060 3244
rect 4492 3176 4500 3184
rect 4764 3176 4772 3184
rect 4876 3176 4884 3184
rect 4460 3156 4468 3164
rect 4604 3156 4612 3164
rect 4716 3156 4724 3164
rect 4508 3136 4516 3144
rect 4412 3116 4420 3124
rect 4444 3076 4452 3084
rect 4412 3056 4420 3064
rect 4428 3056 4436 3064
rect 4396 3016 4404 3024
rect 4412 2936 4420 2944
rect 4428 2936 4436 2944
rect 4460 2956 4468 2964
rect 4444 2916 4452 2924
rect 4460 2916 4468 2924
rect 4396 2896 4404 2904
rect 4444 2896 4452 2904
rect 4412 2716 4420 2724
rect 4476 2896 4484 2904
rect 4636 3136 4644 3144
rect 4684 3136 4692 3144
rect 4524 3116 4532 3124
rect 4572 3116 4580 3124
rect 4540 3076 4548 3084
rect 4524 3056 4532 3064
rect 4556 3056 4564 3064
rect 4540 3036 4548 3044
rect 4540 3016 4548 3024
rect 4540 2956 4548 2964
rect 4652 3116 4660 3124
rect 4636 3056 4644 3064
rect 4636 3036 4644 3044
rect 4668 3036 4676 3044
rect 4588 2956 4596 2964
rect 4556 2936 4564 2944
rect 4732 3116 4740 3124
rect 4700 3076 4708 3084
rect 4812 3096 4820 3104
rect 4956 3096 4964 3104
rect 4988 3096 4996 3104
rect 4732 2936 4740 2944
rect 4620 2916 4628 2924
rect 4508 2896 4516 2904
rect 4604 2896 4612 2904
rect 4700 2896 4708 2904
rect 4572 2836 4580 2844
rect 4684 2836 4692 2844
rect 4540 2796 4548 2804
rect 4748 2816 4756 2824
rect 4668 2756 4676 2764
rect 4764 2756 4772 2764
rect 4508 2736 4516 2744
rect 4620 2736 4628 2744
rect 4684 2736 4692 2744
rect 4492 2696 4500 2704
rect 4460 2676 4468 2684
rect 4268 2616 4276 2624
rect 4316 2616 4324 2624
rect 4204 2576 4212 2584
rect 4300 2576 4308 2584
rect 4156 2556 4164 2564
rect 4188 2556 4196 2564
rect 4188 2516 4196 2524
rect 4108 2496 4116 2504
rect 4108 2456 4116 2464
rect 4076 2376 4084 2384
rect 3916 2356 3924 2364
rect 3852 2216 3860 2224
rect 3788 2156 3796 2164
rect 3836 2156 3844 2164
rect 3820 2116 3828 2124
rect 3756 2016 3764 2024
rect 3756 1996 3764 2004
rect 3708 1956 3716 1964
rect 3756 1956 3764 1964
rect 3724 1936 3732 1944
rect 3836 2096 3844 2104
rect 3820 1956 3828 1964
rect 3900 2096 3908 2104
rect 3852 2076 3860 2084
rect 3788 1916 3796 1924
rect 3596 1896 3604 1904
rect 3612 1896 3620 1904
rect 3692 1896 3700 1904
rect 3788 1896 3796 1904
rect 3836 1896 3844 1904
rect 3836 1876 3844 1884
rect 3820 1856 3828 1864
rect 3644 1796 3652 1804
rect 3740 1796 3748 1804
rect 3772 1796 3780 1804
rect 3628 1776 3636 1784
rect 3500 1756 3508 1764
rect 3532 1736 3540 1744
rect 3580 1736 3588 1744
rect 3596 1736 3604 1744
rect 3500 1676 3508 1684
rect 3516 1636 3524 1644
rect 3660 1756 3668 1764
rect 3900 1956 3908 1964
rect 3868 1916 3876 1924
rect 3964 2276 3972 2284
rect 3948 2116 3956 2124
rect 3996 2296 4004 2304
rect 4060 2296 4068 2304
rect 4092 2296 4100 2304
rect 4044 2156 4052 2164
rect 4060 2156 4068 2164
rect 4140 2376 4148 2384
rect 4268 2476 4276 2484
rect 4348 2456 4356 2464
rect 4476 2616 4484 2624
rect 4956 3076 4964 3084
rect 4924 3056 4932 3064
rect 4940 3036 4948 3044
rect 4908 3016 4916 3024
rect 4972 3056 4980 3064
rect 4972 3016 4980 3024
rect 4860 2936 4868 2944
rect 5068 3096 5076 3104
rect 5068 3036 5076 3044
rect 5164 3136 5172 3144
rect 5132 3116 5140 3124
rect 5116 3096 5124 3104
rect 5116 3076 5124 3084
rect 5228 3276 5236 3284
rect 5292 3316 5300 3324
rect 5260 3176 5268 3184
rect 5324 3176 5332 3184
rect 5196 3116 5204 3124
rect 5404 3416 5412 3424
rect 5436 3396 5444 3404
rect 5484 3456 5492 3464
rect 5468 3436 5476 3444
rect 5436 3356 5444 3364
rect 5404 3316 5412 3324
rect 5516 3456 5524 3464
rect 5500 3416 5508 3424
rect 5676 3656 5684 3664
rect 5548 3636 5556 3644
rect 5580 3636 5588 3644
rect 5548 3496 5556 3504
rect 5612 3516 5620 3524
rect 5644 3516 5652 3524
rect 5580 3456 5588 3464
rect 5692 3476 5700 3484
rect 5676 3436 5684 3444
rect 5660 3416 5668 3424
rect 5580 3376 5588 3384
rect 5612 3376 5620 3384
rect 5596 3356 5604 3364
rect 5500 3336 5508 3344
rect 5548 3336 5556 3344
rect 5500 3316 5508 3324
rect 5788 3716 5796 3724
rect 5852 3736 5860 3744
rect 5788 3696 5796 3704
rect 5820 3696 5828 3704
rect 5836 3696 5844 3704
rect 5740 3676 5748 3684
rect 5788 3656 5796 3664
rect 5788 3556 5796 3564
rect 5724 3536 5732 3544
rect 5772 3516 5780 3524
rect 5804 3536 5812 3544
rect 5756 3496 5764 3504
rect 5852 3516 5860 3524
rect 5772 3456 5780 3464
rect 5820 3456 5828 3464
rect 5708 3376 5716 3384
rect 5660 3316 5668 3324
rect 5564 3276 5572 3284
rect 5708 3356 5716 3364
rect 5740 3276 5748 3284
rect 5852 3416 5860 3424
rect 5788 3316 5796 3324
rect 5788 3256 5796 3264
rect 5820 3276 5828 3284
rect 5932 3796 5940 3804
rect 5916 3716 5924 3724
rect 6060 3856 6068 3864
rect 6060 3836 6068 3844
rect 6350 4206 6358 4214
rect 6364 4206 6372 4214
rect 6378 4206 6386 4214
rect 6268 4156 6276 4164
rect 6316 4156 6324 4164
rect 6252 4136 6260 4144
rect 6492 4256 6500 4264
rect 6588 4256 6596 4264
rect 6460 4196 6468 4204
rect 6556 4216 6564 4224
rect 6492 4176 6500 4184
rect 6524 4176 6532 4184
rect 6620 4236 6628 4244
rect 6652 4216 6660 4224
rect 6572 4196 6580 4204
rect 6652 4196 6660 4204
rect 6780 4216 6788 4224
rect 6668 4156 6676 4164
rect 6684 4156 6692 4164
rect 6476 4136 6484 4144
rect 6508 4116 6516 4124
rect 6620 4096 6628 4104
rect 6348 3996 6356 4004
rect 6428 3976 6436 3984
rect 6268 3956 6276 3964
rect 6540 3956 6548 3964
rect 6236 3916 6244 3924
rect 6220 3896 6228 3904
rect 6076 3796 6084 3804
rect 6140 3796 6148 3804
rect 6012 3756 6020 3764
rect 5980 3736 5988 3744
rect 5948 3676 5956 3684
rect 5964 3676 5972 3684
rect 5916 3656 5924 3664
rect 5900 3536 5908 3544
rect 5932 3596 5940 3604
rect 5916 3516 5924 3524
rect 5900 3496 5908 3504
rect 5964 3616 5972 3624
rect 5980 3596 5988 3604
rect 5996 3516 6004 3524
rect 6028 3716 6036 3724
rect 6044 3716 6052 3724
rect 6108 3716 6116 3724
rect 6124 3676 6132 3684
rect 6044 3616 6052 3624
rect 6028 3596 6036 3604
rect 6060 3516 6068 3524
rect 5980 3476 5988 3484
rect 5900 3416 5908 3424
rect 5884 3376 5892 3384
rect 5900 3336 5908 3344
rect 5884 3296 5892 3304
rect 5356 3116 5364 3124
rect 5404 3116 5412 3124
rect 5484 3116 5492 3124
rect 5852 3116 5860 3124
rect 5196 3076 5204 3084
rect 5340 3076 5348 3084
rect 5932 3256 5940 3264
rect 6060 3456 6068 3464
rect 6044 3436 6052 3444
rect 6060 3376 6068 3384
rect 6092 3536 6100 3544
rect 6124 3536 6132 3544
rect 6092 3456 6100 3464
rect 6076 3356 6084 3364
rect 6124 3436 6132 3444
rect 6012 3336 6020 3344
rect 6076 3336 6084 3344
rect 6028 3256 6036 3264
rect 6028 3236 6036 3244
rect 6124 3276 6132 3284
rect 5948 3216 5956 3224
rect 5964 3216 5972 3224
rect 6108 3216 6116 3224
rect 5932 3136 5940 3144
rect 5676 3096 5684 3104
rect 5708 3096 5716 3104
rect 5756 3096 5764 3104
rect 5916 3096 5924 3104
rect 5084 2936 5092 2944
rect 5148 2936 5156 2944
rect 4796 2896 4804 2904
rect 4908 2896 4916 2904
rect 5164 2916 5172 2924
rect 4814 2806 4822 2814
rect 4828 2806 4836 2814
rect 4842 2806 4850 2814
rect 4796 2776 4804 2784
rect 4668 2716 4676 2724
rect 4716 2716 4724 2724
rect 4780 2716 4788 2724
rect 4892 2716 4900 2724
rect 4556 2696 4564 2704
rect 4748 2696 4756 2704
rect 4556 2676 4564 2684
rect 4636 2676 4644 2684
rect 4732 2676 4740 2684
rect 4556 2656 4564 2664
rect 4588 2656 4596 2664
rect 4652 2656 4660 2664
rect 4556 2636 4564 2644
rect 4620 2636 4628 2644
rect 4604 2596 4612 2604
rect 4652 2616 4660 2624
rect 4460 2576 4468 2584
rect 4540 2576 4548 2584
rect 4604 2576 4612 2584
rect 4444 2556 4452 2564
rect 4380 2516 4388 2524
rect 4396 2516 4404 2524
rect 4396 2476 4404 2484
rect 4364 2436 4372 2444
rect 4316 2416 4324 2424
rect 4300 2376 4308 2384
rect 4252 2356 4260 2364
rect 4428 2456 4436 2464
rect 4428 2436 4436 2444
rect 4236 2336 4244 2344
rect 4332 2336 4340 2344
rect 4396 2336 4404 2344
rect 4268 2316 4276 2324
rect 4364 2296 4372 2304
rect 4412 2296 4420 2304
rect 4380 2236 4388 2244
rect 4124 2136 4132 2144
rect 4092 2116 4100 2124
rect 4028 2096 4036 2104
rect 4060 2096 4068 2104
rect 3980 2056 3988 2064
rect 3980 2036 3988 2044
rect 3964 2016 3972 2024
rect 3932 1996 3940 2004
rect 3948 1956 3956 1964
rect 3884 1876 3892 1884
rect 3916 1876 3924 1884
rect 3916 1836 3924 1844
rect 3852 1796 3860 1804
rect 3932 1796 3940 1804
rect 3756 1756 3764 1764
rect 3804 1756 3812 1764
rect 3820 1756 3828 1764
rect 3676 1736 3684 1744
rect 3852 1736 3860 1744
rect 3788 1696 3796 1704
rect 3820 1696 3828 1704
rect 3900 1736 3908 1744
rect 3740 1656 3748 1664
rect 3868 1656 3876 1664
rect 3948 1656 3956 1664
rect 3580 1636 3588 1644
rect 3676 1616 3684 1624
rect 3564 1596 3572 1604
rect 3596 1556 3604 1564
rect 3532 1516 3540 1524
rect 3708 1596 3716 1604
rect 3628 1476 3636 1484
rect 3692 1476 3700 1484
rect 3548 1436 3556 1444
rect 3532 1356 3540 1364
rect 3516 1336 3524 1344
rect 3116 1276 3124 1284
rect 2796 1216 2804 1224
rect 2796 1196 2804 1204
rect 2828 1116 2836 1124
rect 2732 1096 2740 1104
rect 2812 1096 2820 1104
rect 2716 1076 2724 1084
rect 3276 1276 3284 1284
rect 3148 1176 3156 1184
rect 2876 1156 2884 1164
rect 3068 1156 3076 1164
rect 3404 1136 3412 1144
rect 2940 1102 2948 1104
rect 2940 1096 2948 1102
rect 3084 1076 3092 1084
rect 2668 1056 2676 1064
rect 2844 1056 2852 1064
rect 2908 1056 2916 1064
rect 2636 1036 2644 1044
rect 2780 1036 2788 1044
rect 2812 1036 2820 1044
rect 2716 976 2724 984
rect 2636 956 2644 964
rect 2700 956 2708 964
rect 2716 936 2724 944
rect 2684 916 2692 924
rect 2780 918 2788 924
rect 2780 916 2788 918
rect 2620 836 2628 844
rect 2572 756 2580 764
rect 2540 736 2548 744
rect 2572 736 2580 744
rect 2556 676 2564 684
rect 2604 716 2612 724
rect 2588 696 2596 704
rect 2684 896 2692 904
rect 2748 896 2756 904
rect 2684 736 2692 744
rect 2700 716 2708 724
rect 2412 576 2420 584
rect 2348 556 2356 564
rect 2444 556 2452 564
rect 2476 556 2484 564
rect 2332 536 2340 544
rect 2556 536 2564 544
rect 1980 516 1988 524
rect 2028 516 2036 524
rect 2076 516 2084 524
rect 2252 516 2260 524
rect 1932 476 1940 484
rect 2348 516 2356 524
rect 2444 496 2452 504
rect 2364 476 2372 484
rect 2396 476 2404 484
rect 2028 456 2036 464
rect 1932 316 1940 324
rect 1820 296 1828 304
rect 1900 296 1908 304
rect 2012 296 2020 304
rect 1740 216 1748 224
rect 1756 156 1764 164
rect 1724 136 1732 144
rect 2444 336 2452 344
rect 2620 596 2628 604
rect 2748 696 2756 704
rect 2764 696 2772 704
rect 2668 676 2676 684
rect 2780 676 2788 684
rect 2716 656 2724 664
rect 2668 596 2676 604
rect 2748 596 2756 604
rect 2636 556 2644 564
rect 2748 556 2756 564
rect 2652 536 2660 544
rect 2604 516 2612 524
rect 2684 516 2692 524
rect 2508 496 2516 504
rect 2572 496 2580 504
rect 2684 476 2692 484
rect 2588 356 2596 364
rect 2060 316 2068 324
rect 2380 316 2388 324
rect 2156 296 2164 304
rect 2204 296 2212 304
rect 2396 296 2404 304
rect 2412 296 2420 304
rect 1884 236 1892 244
rect 1868 216 1876 224
rect 1900 176 1908 184
rect 1692 116 1700 124
rect 1852 116 1860 124
rect 1884 116 1892 124
rect 1836 96 1844 104
rect 1996 176 2004 184
rect 2028 176 2036 184
rect 1964 156 1972 164
rect 2236 196 2244 204
rect 2316 196 2324 204
rect 2108 176 2116 184
rect 2172 176 2180 184
rect 2124 156 2132 164
rect 2172 156 2180 164
rect 2188 156 2196 164
rect 2236 156 2244 164
rect 2156 136 2164 144
rect 2668 336 2676 344
rect 2476 316 2484 324
rect 2524 296 2532 304
rect 2540 276 2548 284
rect 2476 256 2484 264
rect 2508 176 2516 184
rect 2556 176 2564 184
rect 2252 136 2260 144
rect 2428 136 2436 144
rect 2524 136 2532 144
rect 2300 116 2308 124
rect 2316 116 2324 124
rect 2956 1036 2964 1044
rect 2908 1016 2916 1024
rect 2908 976 2916 984
rect 2892 956 2900 964
rect 2924 956 2932 964
rect 2844 736 2852 744
rect 2844 716 2852 724
rect 2828 696 2836 704
rect 2844 636 2852 644
rect 2876 596 2884 604
rect 2812 556 2820 564
rect 2844 536 2852 544
rect 2732 516 2740 524
rect 2796 516 2804 524
rect 3052 976 3060 984
rect 3004 936 3012 944
rect 2972 916 2980 924
rect 3068 956 3076 964
rect 2908 856 2916 864
rect 3068 856 3076 864
rect 3244 1096 3252 1104
rect 3292 1096 3300 1104
rect 3388 1096 3396 1104
rect 3436 1096 3444 1104
rect 3212 1056 3220 1064
rect 3116 976 3124 984
rect 3228 976 3236 984
rect 3180 956 3188 964
rect 3228 956 3236 964
rect 3132 936 3140 944
rect 3196 936 3204 944
rect 3228 936 3236 944
rect 3276 1076 3284 1084
rect 3372 1076 3380 1084
rect 3278 1006 3286 1014
rect 3292 1006 3300 1014
rect 3306 1006 3314 1014
rect 3244 916 3252 924
rect 3260 896 3268 904
rect 3356 1036 3364 1044
rect 3356 916 3364 924
rect 3500 1276 3508 1284
rect 3596 1456 3604 1464
rect 3932 1636 3940 1644
rect 3724 1536 3732 1544
rect 3932 1536 3940 1544
rect 4012 1936 4020 1944
rect 3996 1916 4004 1924
rect 3996 1816 4004 1824
rect 4044 1916 4052 1924
rect 4028 1896 4036 1904
rect 4076 1956 4084 1964
rect 4060 1856 4068 1864
rect 4172 2156 4180 2164
rect 4156 1996 4164 2004
rect 4140 1976 4148 1984
rect 4108 1896 4116 1904
rect 4236 2136 4244 2144
rect 4284 2136 4292 2144
rect 4348 2216 4356 2224
rect 4412 2216 4420 2224
rect 4236 2056 4244 2064
rect 4188 1916 4196 1924
rect 4284 1976 4292 1984
rect 4172 1896 4180 1904
rect 4220 1896 4228 1904
rect 4108 1876 4116 1884
rect 4076 1816 4084 1824
rect 4060 1796 4068 1804
rect 4316 1936 4324 1944
rect 4124 1776 4132 1784
rect 4268 1796 4276 1804
rect 4412 2136 4420 2144
rect 4540 2556 4548 2564
rect 4572 2556 4580 2564
rect 4476 2516 4484 2524
rect 4540 2516 4548 2524
rect 4556 2496 4564 2504
rect 4476 2476 4484 2484
rect 4444 2296 4452 2304
rect 4508 2376 4516 2384
rect 4588 2416 4596 2424
rect 4588 2396 4596 2404
rect 4556 2336 4564 2344
rect 4492 2316 4500 2324
rect 4524 2316 4532 2324
rect 4572 2316 4580 2324
rect 4460 2236 4468 2244
rect 4508 2256 4516 2264
rect 4540 2256 4548 2264
rect 4492 2216 4500 2224
rect 4476 2196 4484 2204
rect 4492 2176 4500 2184
rect 4444 2156 4452 2164
rect 4476 2156 4484 2164
rect 4380 2116 4388 2124
rect 4524 2236 4532 2244
rect 4636 2556 4644 2564
rect 4748 2556 4756 2564
rect 4684 2536 4692 2544
rect 4748 2536 4756 2544
rect 4620 2476 4628 2484
rect 4668 2336 4676 2344
rect 4636 2316 4644 2324
rect 4780 2596 4788 2604
rect 4828 2596 4836 2604
rect 4764 2476 4772 2484
rect 4764 2456 4772 2464
rect 4716 2396 4724 2404
rect 4700 2316 4708 2324
rect 4748 2296 4756 2304
rect 4814 2406 4822 2414
rect 4828 2406 4836 2414
rect 4842 2406 4850 2414
rect 4812 2376 4820 2384
rect 4780 2316 4788 2324
rect 4652 2256 4660 2264
rect 4684 2256 4692 2264
rect 4780 2256 4788 2264
rect 4556 2236 4564 2244
rect 4572 2216 4580 2224
rect 4652 2216 4660 2224
rect 4588 2196 4596 2204
rect 4636 2016 4644 2024
rect 4508 1916 4516 1924
rect 4588 1916 4596 1924
rect 4396 1896 4404 1904
rect 4364 1856 4372 1864
rect 4396 1796 4404 1804
rect 4252 1776 4260 1784
rect 4348 1776 4356 1784
rect 4108 1736 4116 1744
rect 4140 1736 4148 1744
rect 4316 1756 4324 1764
rect 4380 1756 4388 1764
rect 4364 1736 4372 1744
rect 4028 1716 4036 1724
rect 4012 1676 4020 1684
rect 3980 1556 3988 1564
rect 4444 1796 4452 1804
rect 4412 1736 4420 1744
rect 4716 2196 4724 2204
rect 4876 2356 4884 2364
rect 4828 2316 4836 2324
rect 4828 2296 4836 2304
rect 4844 2236 4852 2244
rect 4892 2236 4900 2244
rect 4796 2156 4804 2164
rect 4668 2116 4676 2124
rect 4716 1936 4724 1944
rect 4814 2006 4822 2014
rect 4828 2006 4836 2014
rect 4842 2006 4850 2014
rect 4876 1936 4884 1944
rect 4892 1936 4900 1944
rect 4780 1896 4788 1904
rect 4812 1896 4820 1904
rect 4860 1896 4868 1904
rect 4492 1856 4500 1864
rect 4620 1856 4628 1864
rect 4524 1836 4532 1844
rect 4476 1796 4484 1804
rect 4460 1756 4468 1764
rect 4444 1716 4452 1724
rect 4556 1836 4564 1844
rect 4540 1816 4548 1824
rect 4492 1696 4500 1704
rect 4188 1676 4196 1684
rect 4076 1636 4084 1644
rect 4444 1676 4452 1684
rect 4812 1856 4820 1864
rect 4764 1836 4772 1844
rect 4780 1836 4788 1844
rect 4684 1816 4692 1824
rect 4652 1796 4660 1804
rect 4636 1756 4644 1764
rect 4700 1756 4708 1764
rect 4620 1716 4628 1724
rect 4668 1716 4676 1724
rect 4076 1596 4084 1604
rect 4092 1596 4100 1604
rect 4412 1596 4420 1604
rect 4044 1556 4052 1564
rect 4252 1556 4260 1564
rect 4204 1536 4212 1544
rect 4044 1516 4052 1524
rect 4140 1516 4148 1524
rect 4172 1516 4180 1524
rect 4316 1516 4324 1524
rect 4428 1516 4436 1524
rect 3852 1496 3860 1504
rect 3964 1496 3972 1504
rect 3596 1376 3604 1384
rect 3628 1316 3636 1324
rect 3484 1076 3492 1084
rect 3468 1036 3476 1044
rect 3452 976 3460 984
rect 3564 1196 3572 1204
rect 3564 1176 3572 1184
rect 3596 1176 3604 1184
rect 3548 1136 3556 1144
rect 3692 1136 3700 1144
rect 3532 1056 3540 1064
rect 3612 1056 3620 1064
rect 3564 1036 3572 1044
rect 3660 1096 3668 1104
rect 3724 1376 3732 1384
rect 3740 1316 3748 1324
rect 3740 1296 3748 1304
rect 3756 1176 3764 1184
rect 3916 1476 3924 1484
rect 3884 1456 3892 1464
rect 3836 1416 3844 1424
rect 3804 1396 3812 1404
rect 3980 1456 3988 1464
rect 4156 1496 4164 1504
rect 4060 1456 4068 1464
rect 4076 1456 4084 1464
rect 4108 1456 4116 1464
rect 4076 1416 4084 1424
rect 4092 1416 4100 1424
rect 4108 1416 4116 1424
rect 3820 1376 3828 1384
rect 4076 1376 4084 1384
rect 3868 1356 3876 1364
rect 3900 1356 3908 1364
rect 3788 1216 3796 1224
rect 3708 1096 3716 1104
rect 3660 1076 3668 1084
rect 3692 1076 3700 1084
rect 3724 1080 3732 1084
rect 3724 1076 3732 1080
rect 3708 1036 3716 1044
rect 3692 956 3700 964
rect 3708 936 3716 944
rect 3500 916 3508 924
rect 3548 916 3556 924
rect 3596 916 3604 924
rect 3436 896 3444 904
rect 3404 856 3412 864
rect 3180 816 3188 824
rect 3004 736 3012 744
rect 3052 736 3060 744
rect 2924 716 2932 724
rect 2940 696 2948 704
rect 2924 676 2932 684
rect 3036 676 3044 684
rect 3084 776 3092 784
rect 3132 776 3140 784
rect 3340 736 3348 744
rect 3372 816 3380 824
rect 3660 916 3668 924
rect 3644 856 3652 864
rect 3676 856 3684 864
rect 3660 776 3668 784
rect 3628 716 3636 724
rect 3340 696 3348 704
rect 3516 702 3524 704
rect 3516 696 3524 702
rect 3260 676 3268 684
rect 3484 676 3492 684
rect 3132 656 3140 664
rect 3452 656 3460 664
rect 3244 636 3252 644
rect 3132 556 3140 564
rect 2924 516 2932 524
rect 3084 516 3092 524
rect 2956 496 2964 504
rect 2988 436 2996 444
rect 2892 416 2900 424
rect 2844 376 2852 384
rect 2812 356 2820 364
rect 2828 356 2836 364
rect 2748 316 2756 324
rect 2716 296 2724 304
rect 2700 276 2708 284
rect 2620 256 2628 264
rect 2620 196 2628 204
rect 2732 256 2740 264
rect 2636 156 2644 164
rect 2812 296 2820 304
rect 2908 376 2916 384
rect 2956 376 2964 384
rect 2908 336 2916 344
rect 2956 336 2964 344
rect 2860 316 2868 324
rect 2828 276 2836 284
rect 2876 276 2884 284
rect 2764 256 2772 264
rect 2828 256 2836 264
rect 2748 176 2756 184
rect 2796 176 2804 184
rect 2764 156 2772 164
rect 2732 136 2740 144
rect 2748 136 2756 144
rect 2780 116 2788 124
rect 3052 396 3060 404
rect 3020 356 3028 364
rect 2988 296 2996 304
rect 3100 376 3108 384
rect 3116 376 3124 384
rect 3180 316 3188 324
rect 3132 276 3140 284
rect 3068 256 3076 264
rect 3164 236 3172 244
rect 2924 176 2932 184
rect 2956 176 2964 184
rect 3004 176 3012 184
rect 3036 176 3044 184
rect 2892 156 2900 164
rect 2908 136 2916 144
rect 2844 116 2852 124
rect 2908 116 2916 124
rect 3278 606 3286 614
rect 3292 606 3300 614
rect 3306 606 3314 614
rect 3436 576 3444 584
rect 3644 596 3652 604
rect 3644 576 3652 584
rect 3340 536 3348 544
rect 3516 536 3524 544
rect 3516 516 3524 524
rect 3260 436 3268 444
rect 3436 436 3444 444
rect 3340 356 3348 364
rect 3292 316 3300 324
rect 3356 336 3364 344
rect 3388 316 3396 324
rect 3420 296 3428 304
rect 3404 276 3412 284
rect 3278 206 3286 214
rect 3292 206 3300 214
rect 3306 206 3314 214
rect 3388 176 3396 184
rect 3020 156 3028 164
rect 3228 156 3236 164
rect 3660 416 3668 424
rect 3644 376 3652 384
rect 3692 696 3700 704
rect 3708 656 3716 664
rect 3740 1016 3748 1024
rect 3740 956 3748 964
rect 3772 1136 3780 1144
rect 4012 1336 4020 1344
rect 4124 1336 4132 1344
rect 3964 1316 3972 1324
rect 4060 1316 4068 1324
rect 3980 1296 3988 1304
rect 3884 1276 3892 1284
rect 3932 1276 3940 1284
rect 4044 1276 4052 1284
rect 3884 1156 3892 1164
rect 4092 1156 4100 1164
rect 4012 1116 4020 1124
rect 4044 1116 4052 1124
rect 3964 1096 3972 1104
rect 3980 1096 3988 1104
rect 3868 1076 3876 1084
rect 3884 1056 3892 1064
rect 3836 1036 3844 1044
rect 4076 1080 4084 1084
rect 4076 1076 4084 1080
rect 4028 1056 4036 1064
rect 4076 1056 4084 1064
rect 3964 1016 3972 1024
rect 3932 996 3940 1004
rect 3932 976 3940 984
rect 3948 976 3956 984
rect 3804 956 3812 964
rect 3756 936 3764 944
rect 3788 936 3796 944
rect 3852 936 3860 944
rect 3916 916 3924 924
rect 3980 976 3988 984
rect 3964 916 3972 924
rect 3916 896 3924 904
rect 3836 876 3844 884
rect 3884 876 3892 884
rect 3900 876 3908 884
rect 3868 856 3876 864
rect 3788 756 3796 764
rect 3852 716 3860 724
rect 3964 796 3972 804
rect 3900 716 3908 724
rect 3756 676 3764 684
rect 3740 656 3748 664
rect 3932 696 3940 704
rect 3804 676 3812 684
rect 4284 1496 4292 1504
rect 4364 1496 4372 1504
rect 4380 1496 4388 1504
rect 4396 1496 4404 1504
rect 4188 1476 4196 1484
rect 4204 1476 4212 1484
rect 4316 1476 4324 1484
rect 4204 1396 4212 1404
rect 4172 1316 4180 1324
rect 4188 1316 4196 1324
rect 4204 1296 4212 1304
rect 4300 1416 4308 1424
rect 4364 1476 4372 1484
rect 4348 1376 4356 1384
rect 4348 1336 4356 1344
rect 4396 1476 4404 1484
rect 4492 1496 4500 1504
rect 4524 1502 4532 1504
rect 4524 1496 4532 1502
rect 4444 1476 4452 1484
rect 4428 1456 4436 1464
rect 4460 1416 4468 1424
rect 4428 1396 4436 1404
rect 4332 1316 4340 1324
rect 4364 1316 4372 1324
rect 4268 1276 4276 1284
rect 4316 1276 4324 1284
rect 4236 1256 4244 1264
rect 4284 1256 4292 1264
rect 4236 1216 4244 1224
rect 4188 1176 4196 1184
rect 4220 1176 4228 1184
rect 4140 1096 4148 1104
rect 4140 1076 4148 1084
rect 4156 1076 4164 1084
rect 4124 956 4132 964
rect 4044 916 4052 924
rect 4044 876 4052 884
rect 3996 856 4004 864
rect 4028 856 4036 864
rect 4012 696 4020 704
rect 4028 696 4036 704
rect 4140 936 4148 944
rect 4204 1056 4212 1064
rect 4188 1016 4196 1024
rect 4252 1096 4260 1104
rect 4268 1076 4276 1084
rect 4236 1036 4244 1044
rect 4268 1016 4276 1024
rect 4220 976 4228 984
rect 4268 956 4276 964
rect 4156 916 4164 924
rect 4108 896 4116 904
rect 4092 876 4100 884
rect 4108 816 4116 824
rect 4108 796 4116 804
rect 4380 1256 4388 1264
rect 4492 1396 4500 1404
rect 4460 1316 4468 1324
rect 4460 1296 4468 1304
rect 4524 1316 4532 1324
rect 4492 1256 4500 1264
rect 4348 1102 4356 1104
rect 4348 1096 4356 1102
rect 4348 1056 4356 1064
rect 4524 1096 4532 1104
rect 4460 1036 4468 1044
rect 4476 1016 4484 1024
rect 4508 1016 4516 1024
rect 4412 976 4420 984
rect 4476 976 4484 984
rect 4380 956 4388 964
rect 4428 956 4436 964
rect 4460 956 4468 964
rect 4300 936 4308 944
rect 4204 876 4212 884
rect 4380 916 4388 924
rect 4268 776 4276 784
rect 4236 736 4244 744
rect 4156 716 4164 724
rect 4092 696 4100 704
rect 4108 696 4116 704
rect 4140 696 4148 704
rect 4076 676 4084 684
rect 4188 676 4196 684
rect 3820 656 3828 664
rect 3788 636 3796 644
rect 3724 576 3732 584
rect 3708 516 3716 524
rect 3724 496 3732 504
rect 3932 576 3940 584
rect 4028 616 4036 624
rect 4220 596 4228 604
rect 4124 576 4132 584
rect 4300 796 4308 804
rect 4300 676 4308 684
rect 4284 656 4292 664
rect 4268 576 4276 584
rect 4252 556 4260 564
rect 4028 536 4036 544
rect 3868 518 3876 524
rect 3868 516 3876 518
rect 3948 516 3956 524
rect 4060 518 4068 524
rect 4060 516 4068 518
rect 4188 516 4196 524
rect 3852 496 3860 504
rect 3804 476 3812 484
rect 4124 476 4132 484
rect 4172 476 4180 484
rect 3772 456 3780 464
rect 3756 396 3764 404
rect 3548 336 3556 344
rect 3484 316 3492 324
rect 3596 316 3604 324
rect 3484 296 3492 304
rect 3548 296 3556 304
rect 3484 276 3492 284
rect 3532 276 3540 284
rect 3756 376 3764 384
rect 3676 356 3684 364
rect 3692 336 3700 344
rect 3628 256 3636 264
rect 3676 256 3684 264
rect 3532 236 3540 244
rect 3724 296 3732 304
rect 3948 436 3956 444
rect 3804 356 3812 364
rect 3916 336 3924 344
rect 3900 316 3908 324
rect 3932 316 3940 324
rect 3884 296 3892 304
rect 3900 296 3908 304
rect 3708 256 3716 264
rect 3772 256 3780 264
rect 3820 256 3828 264
rect 3420 176 3428 184
rect 3708 216 3716 224
rect 3724 176 3732 184
rect 2988 136 2996 144
rect 3132 136 3140 144
rect 3308 136 3316 144
rect 3436 136 3444 144
rect 3532 136 3540 144
rect 3004 116 3012 124
rect 3340 116 3348 124
rect 3452 116 3460 124
rect 3884 256 3892 264
rect 3916 256 3924 264
rect 3932 256 3940 264
rect 3820 236 3828 244
rect 3868 236 3876 244
rect 3836 216 3844 224
rect 3772 156 3780 164
rect 3740 136 3748 144
rect 3788 136 3796 144
rect 3820 136 3828 144
rect 3852 156 3860 164
rect 3916 216 3924 224
rect 4028 356 4036 364
rect 3964 336 3972 344
rect 4108 302 4116 304
rect 4108 296 4116 302
rect 3996 276 4004 284
rect 3980 256 3988 264
rect 3660 116 3668 124
rect 3692 116 3700 124
rect 3820 116 3828 124
rect 3900 116 3908 124
rect 3948 116 3956 124
rect 1900 96 1908 104
rect 1916 96 1924 104
rect 1948 96 1956 104
rect 1980 96 1988 104
rect 1996 96 2004 104
rect 2044 96 2052 104
rect 2460 96 2468 104
rect 2572 96 2580 104
rect 2604 96 2612 104
rect 2668 96 2676 104
rect 3468 96 3476 104
rect 140 76 148 84
rect 204 76 212 84
rect 764 76 772 84
rect 940 76 948 84
rect 1388 76 1396 84
rect 1532 76 1540 84
rect 1564 76 1572 84
rect 1756 76 1764 84
rect 1868 76 1876 84
rect 1884 76 1892 84
rect 4204 456 4212 464
rect 4236 336 4244 344
rect 4508 916 4516 924
rect 4652 1576 4660 1584
rect 4716 1716 4724 1724
rect 4700 1536 4708 1544
rect 4588 1516 4596 1524
rect 4956 2856 4964 2864
rect 5068 2896 5076 2904
rect 5004 2716 5012 2724
rect 5004 2696 5012 2704
rect 4956 2556 4964 2564
rect 5004 2556 5012 2564
rect 5660 3076 5668 3084
rect 5564 3056 5572 3064
rect 5532 3036 5540 3044
rect 5564 3036 5572 3044
rect 5260 2976 5268 2984
rect 5388 2976 5396 2984
rect 5356 2936 5364 2944
rect 5212 2876 5220 2884
rect 5196 2856 5204 2864
rect 5308 2856 5316 2864
rect 5068 2756 5076 2764
rect 5084 2716 5092 2724
rect 5020 2516 5028 2524
rect 5004 2376 5012 2384
rect 4940 2336 4948 2344
rect 5020 2316 5028 2324
rect 4988 2296 4996 2304
rect 4924 2256 4932 2264
rect 5020 2256 5028 2264
rect 4956 2236 4964 2244
rect 4972 2196 4980 2204
rect 5052 2456 5060 2464
rect 5052 2396 5060 2404
rect 5068 2316 5076 2324
rect 5276 2816 5284 2824
rect 5244 2796 5252 2804
rect 5164 2716 5172 2724
rect 5148 2696 5156 2704
rect 5180 2696 5188 2704
rect 5260 2696 5268 2704
rect 5132 2676 5140 2684
rect 5212 2676 5220 2684
rect 5180 2636 5188 2644
rect 5164 2616 5172 2624
rect 5260 2656 5268 2664
rect 5116 2576 5124 2584
rect 5180 2536 5188 2544
rect 5260 2536 5268 2544
rect 5292 2796 5300 2804
rect 5356 2736 5364 2744
rect 5324 2716 5332 2724
rect 5484 2996 5492 3004
rect 5468 2976 5476 2984
rect 5532 2956 5540 2964
rect 5436 2916 5444 2924
rect 5436 2876 5444 2884
rect 5388 2716 5396 2724
rect 5452 2836 5460 2844
rect 5404 2676 5412 2684
rect 5308 2576 5316 2584
rect 5212 2516 5220 2524
rect 5436 2656 5444 2664
rect 5324 2556 5332 2564
rect 5356 2536 5364 2544
rect 5548 2936 5556 2944
rect 5516 2816 5524 2824
rect 5500 2796 5508 2804
rect 5516 2756 5524 2764
rect 5516 2736 5524 2744
rect 5484 2716 5492 2724
rect 5516 2716 5524 2724
rect 5468 2696 5476 2704
rect 5596 2996 5604 3004
rect 5660 2996 5668 3004
rect 5612 2956 5620 2964
rect 5580 2916 5588 2924
rect 5580 2816 5588 2824
rect 5596 2796 5604 2804
rect 5580 2716 5588 2724
rect 5532 2676 5540 2684
rect 5564 2676 5572 2684
rect 5484 2536 5492 2544
rect 5404 2516 5412 2524
rect 5500 2516 5508 2524
rect 5132 2396 5140 2404
rect 5212 2396 5220 2404
rect 5388 2356 5396 2364
rect 5084 2296 5092 2304
rect 5100 2296 5108 2304
rect 5244 2296 5252 2304
rect 5260 2276 5268 2284
rect 5084 2216 5092 2224
rect 4988 2136 4996 2144
rect 5036 2136 5044 2144
rect 4956 2118 4964 2124
rect 4956 2116 4964 2118
rect 5068 2116 5076 2124
rect 4956 2076 4964 2084
rect 5020 2076 5028 2084
rect 5052 2076 5060 2084
rect 5260 2196 5268 2204
rect 5116 2176 5124 2184
rect 5100 2156 5108 2164
rect 5100 2136 5108 2144
rect 5052 1936 5060 1944
rect 4956 1896 4964 1904
rect 5004 1896 5012 1904
rect 5084 1896 5092 1904
rect 4988 1816 4996 1824
rect 5036 1816 5044 1824
rect 5004 1776 5012 1784
rect 5020 1776 5028 1784
rect 4988 1756 4996 1764
rect 4828 1676 4836 1684
rect 4924 1676 4932 1684
rect 4814 1606 4822 1614
rect 4828 1606 4836 1614
rect 4842 1606 4850 1614
rect 4988 1576 4996 1584
rect 4892 1536 4900 1544
rect 4748 1516 4756 1524
rect 4700 1496 4708 1504
rect 4716 1496 4724 1504
rect 4732 1496 4740 1504
rect 4892 1496 4900 1504
rect 4940 1496 4948 1504
rect 4556 1276 4564 1284
rect 4716 1476 4724 1484
rect 4764 1476 4772 1484
rect 4620 1456 4628 1464
rect 4604 1416 4612 1424
rect 4668 1396 4676 1404
rect 4732 1396 4740 1404
rect 4716 1376 4724 1384
rect 4604 996 4612 1004
rect 4604 956 4612 964
rect 4588 936 4596 944
rect 4556 896 4564 904
rect 4540 876 4548 884
rect 4876 1476 4884 1484
rect 4972 1476 4980 1484
rect 4988 1456 4996 1464
rect 4812 1416 4820 1424
rect 4780 1376 4788 1384
rect 4716 1316 4724 1324
rect 4908 1336 4916 1344
rect 5052 1796 5060 1804
rect 5084 1776 5092 1784
rect 5068 1756 5076 1764
rect 5084 1736 5092 1744
rect 5036 1716 5044 1724
rect 5036 1576 5044 1584
rect 5180 2136 5188 2144
rect 5340 2176 5348 2184
rect 5308 2156 5316 2164
rect 5276 2116 5284 2124
rect 5180 2076 5188 2084
rect 5452 2376 5460 2384
rect 5516 2356 5524 2364
rect 5500 2316 5508 2324
rect 5404 2296 5412 2304
rect 5388 2156 5396 2164
rect 5548 2656 5556 2664
rect 5564 2596 5572 2604
rect 5580 2556 5588 2564
rect 5660 2876 5668 2884
rect 5724 3056 5732 3064
rect 5708 2936 5716 2944
rect 5676 2836 5684 2844
rect 5756 2936 5764 2944
rect 5740 2916 5748 2924
rect 5724 2816 5732 2824
rect 5708 2796 5716 2804
rect 5692 2756 5700 2764
rect 5756 2836 5764 2844
rect 5692 2736 5700 2744
rect 5740 2736 5748 2744
rect 5836 3036 5844 3044
rect 5804 2996 5812 3004
rect 5836 2996 5844 3004
rect 5788 2936 5796 2944
rect 5820 2916 5828 2924
rect 5900 3076 5908 3084
rect 5948 3036 5956 3044
rect 5900 2936 5908 2944
rect 5932 2736 5940 2744
rect 5884 2716 5892 2724
rect 5708 2696 5716 2704
rect 5852 2696 5860 2704
rect 5900 2696 5908 2704
rect 5756 2676 5764 2684
rect 5772 2676 5780 2684
rect 5820 2676 5828 2684
rect 5724 2656 5732 2664
rect 5740 2656 5748 2664
rect 5692 2636 5700 2644
rect 5724 2636 5732 2644
rect 5612 2616 5620 2624
rect 5708 2616 5716 2624
rect 5660 2576 5668 2584
rect 6124 3136 6132 3144
rect 6156 3736 6164 3744
rect 6156 3716 6164 3724
rect 6172 3576 6180 3584
rect 6396 3902 6404 3904
rect 6396 3896 6404 3902
rect 6492 3896 6500 3904
rect 6364 3856 6372 3864
rect 6350 3806 6358 3814
rect 6364 3806 6372 3814
rect 6378 3806 6386 3814
rect 6556 3916 6564 3924
rect 6300 3736 6308 3744
rect 6412 3736 6420 3744
rect 6428 3736 6436 3744
rect 6508 3736 6516 3744
rect 6444 3716 6452 3724
rect 6316 3696 6324 3704
rect 6284 3676 6292 3684
rect 6252 3656 6260 3664
rect 6236 3616 6244 3624
rect 6204 3536 6212 3544
rect 6188 3516 6196 3524
rect 6252 3556 6260 3564
rect 6284 3596 6292 3604
rect 6284 3556 6292 3564
rect 6380 3536 6388 3544
rect 6300 3516 6308 3524
rect 6332 3516 6340 3524
rect 6236 3496 6244 3504
rect 6268 3496 6276 3504
rect 6364 3496 6372 3504
rect 6156 3456 6164 3464
rect 6236 3456 6244 3464
rect 6332 3456 6340 3464
rect 6140 3116 6148 3124
rect 6188 3416 6196 3424
rect 6172 3196 6180 3204
rect 6012 3096 6020 3104
rect 6076 3102 6084 3104
rect 6076 3096 6084 3102
rect 6172 3096 6180 3104
rect 6156 3076 6164 3084
rect 6012 3036 6020 3044
rect 5996 2996 6004 3004
rect 5884 2676 5892 2684
rect 5948 2676 5956 2684
rect 5964 2676 5972 2684
rect 5868 2656 5876 2664
rect 5804 2636 5812 2644
rect 5740 2556 5748 2564
rect 5756 2556 5764 2564
rect 5644 2536 5652 2544
rect 5724 2536 5732 2544
rect 5916 2616 5924 2624
rect 5868 2556 5876 2564
rect 5996 2676 6004 2684
rect 6140 3036 6148 3044
rect 6350 3406 6358 3414
rect 6364 3406 6372 3414
rect 6378 3406 6386 3414
rect 6396 3356 6404 3364
rect 6332 3316 6340 3324
rect 6300 3296 6308 3304
rect 6364 3296 6372 3304
rect 6236 3216 6244 3224
rect 6268 3196 6276 3204
rect 6236 3116 6244 3124
rect 6220 3076 6228 3084
rect 6444 3496 6452 3504
rect 6492 3716 6500 3724
rect 6476 3516 6484 3524
rect 6588 3896 6596 3904
rect 6620 3896 6628 3904
rect 6620 3876 6628 3884
rect 6572 3816 6580 3824
rect 6636 3816 6644 3824
rect 6636 3716 6644 3724
rect 6588 3696 6596 3704
rect 6524 3676 6532 3684
rect 6572 3676 6580 3684
rect 6620 3656 6628 3664
rect 6668 4096 6676 4104
rect 6700 4096 6708 4104
rect 6716 4056 6724 4064
rect 6668 3996 6676 4004
rect 6748 4116 6756 4124
rect 6844 4496 6852 4504
rect 6860 4496 6868 4504
rect 6860 4316 6868 4324
rect 6844 4296 6852 4304
rect 6908 4296 6916 4304
rect 6828 4276 6836 4284
rect 6892 4276 6900 4284
rect 6924 4216 6932 4224
rect 6844 4156 6852 4164
rect 6812 4116 6820 4124
rect 6748 4096 6756 4104
rect 6844 4056 6852 4064
rect 6828 4036 6836 4044
rect 6732 3956 6740 3964
rect 6860 3936 6868 3944
rect 6876 3916 6884 3924
rect 6668 3896 6676 3904
rect 6732 3896 6740 3904
rect 6860 3896 6868 3904
rect 6716 3876 6724 3884
rect 6796 3876 6804 3884
rect 6684 3796 6692 3804
rect 6972 4518 6980 4524
rect 6972 4516 6980 4518
rect 7100 4476 7108 4484
rect 7052 4436 7060 4444
rect 6956 4336 6964 4344
rect 6972 4196 6980 4204
rect 7196 4556 7204 4564
rect 7436 4576 7444 4584
rect 7276 4556 7284 4564
rect 7356 4556 7364 4564
rect 7404 4556 7412 4564
rect 7164 4536 7172 4544
rect 7164 4516 7172 4524
rect 7132 4436 7140 4444
rect 7148 4436 7156 4444
rect 7228 4518 7236 4524
rect 7228 4516 7236 4518
rect 7372 4536 7380 4544
rect 7276 4496 7284 4504
rect 7372 4496 7380 4504
rect 7148 4416 7156 4424
rect 7196 4416 7204 4424
rect 7116 4336 7124 4344
rect 7116 4316 7124 4324
rect 7196 4336 7204 4344
rect 7292 4336 7300 4344
rect 7244 4316 7252 4324
rect 7260 4316 7268 4324
rect 7196 4296 7204 4304
rect 7116 4256 7124 4264
rect 7084 4216 7092 4224
rect 7276 4296 7284 4304
rect 7228 4276 7236 4284
rect 7260 4276 7268 4284
rect 7212 4256 7220 4264
rect 7228 4256 7236 4264
rect 7148 4236 7156 4244
rect 7260 4216 7268 4224
rect 7100 4176 7108 4184
rect 7324 4316 7332 4324
rect 7356 4316 7364 4324
rect 7388 4316 7396 4324
rect 7372 4296 7380 4304
rect 7308 4276 7316 4284
rect 7308 4176 7316 4184
rect 7308 4156 7316 4164
rect 6988 4136 6996 4144
rect 7100 4136 7108 4144
rect 7100 4116 7108 4124
rect 6972 4076 6980 4084
rect 6908 3916 6916 3924
rect 7084 3916 7092 3924
rect 6908 3896 6916 3904
rect 6892 3876 6900 3884
rect 6908 3836 6916 3844
rect 6748 3736 6756 3744
rect 6876 3736 6884 3744
rect 6732 3716 6740 3724
rect 6684 3676 6692 3684
rect 6652 3616 6660 3624
rect 6524 3576 6532 3584
rect 6524 3536 6532 3544
rect 6620 3536 6628 3544
rect 6700 3536 6708 3544
rect 6508 3516 6516 3524
rect 6604 3516 6612 3524
rect 6524 3496 6532 3504
rect 6604 3496 6612 3504
rect 6540 3476 6548 3484
rect 6492 3456 6500 3464
rect 6524 3436 6532 3444
rect 6444 3376 6452 3384
rect 6716 3496 6724 3504
rect 6700 3456 6708 3464
rect 6572 3436 6580 3444
rect 6668 3416 6676 3424
rect 6588 3376 6596 3384
rect 6652 3376 6660 3384
rect 6700 3356 6708 3364
rect 6748 3356 6756 3364
rect 6540 3336 6548 3344
rect 6652 3336 6660 3344
rect 6812 3716 6820 3724
rect 6860 3716 6868 3724
rect 6940 3716 6948 3724
rect 6828 3656 6836 3664
rect 6892 3696 6900 3704
rect 6908 3556 6916 3564
rect 6828 3496 6836 3504
rect 6796 3436 6804 3444
rect 6780 3376 6788 3384
rect 6764 3316 6772 3324
rect 6556 3216 6564 3224
rect 6508 3196 6516 3204
rect 6412 3156 6420 3164
rect 6444 3156 6452 3164
rect 6316 3136 6324 3144
rect 6316 3096 6324 3104
rect 6396 3096 6404 3104
rect 6428 3096 6436 3104
rect 6268 3076 6276 3084
rect 6092 2916 6100 2924
rect 6252 2896 6260 2904
rect 6108 2736 6116 2744
rect 6172 2736 6180 2744
rect 6092 2696 6100 2704
rect 5980 2656 5988 2664
rect 6012 2656 6020 2664
rect 6140 2656 6148 2664
rect 6140 2636 6148 2644
rect 6060 2596 6068 2604
rect 6012 2556 6020 2564
rect 5852 2536 5860 2544
rect 5612 2516 5620 2524
rect 5660 2516 5668 2524
rect 5692 2516 5700 2524
rect 5740 2516 5748 2524
rect 5852 2516 5860 2524
rect 5964 2536 5972 2544
rect 6028 2536 6036 2544
rect 6124 2576 6132 2584
rect 6156 2556 6164 2564
rect 6108 2516 6116 2524
rect 6172 2516 6180 2524
rect 5932 2496 5940 2504
rect 5980 2496 5988 2504
rect 6028 2496 6036 2504
rect 6076 2496 6084 2504
rect 5884 2456 5892 2464
rect 5916 2456 5924 2464
rect 5756 2376 5764 2384
rect 5740 2356 5748 2364
rect 5644 2336 5652 2344
rect 5628 2316 5636 2324
rect 5596 2296 5604 2304
rect 5452 2276 5460 2284
rect 5516 2276 5524 2284
rect 5532 2276 5540 2284
rect 5580 2280 5588 2284
rect 5580 2276 5588 2280
rect 5596 2256 5604 2264
rect 5484 2196 5492 2204
rect 5516 2176 5524 2184
rect 5468 2136 5476 2144
rect 5372 2116 5380 2124
rect 5308 1996 5316 2004
rect 5116 1916 5124 1924
rect 5148 1916 5156 1924
rect 5132 1896 5140 1904
rect 5228 1896 5236 1904
rect 5276 1896 5284 1904
rect 5196 1836 5204 1844
rect 5212 1816 5220 1824
rect 5116 1796 5124 1804
rect 5196 1736 5204 1744
rect 5116 1516 5124 1524
rect 5100 1476 5108 1484
rect 5020 1416 5028 1424
rect 4940 1336 4948 1344
rect 4876 1316 4884 1324
rect 4908 1316 4916 1324
rect 4780 1296 4788 1304
rect 4748 1156 4756 1164
rect 4652 1116 4660 1124
rect 4732 1116 4740 1124
rect 4764 1116 4772 1124
rect 4716 1076 4724 1084
rect 4732 1056 4740 1064
rect 4700 996 4708 1004
rect 4764 1076 4772 1084
rect 4748 1036 4756 1044
rect 4764 996 4772 1004
rect 4684 916 4692 924
rect 4748 896 4756 904
rect 4620 856 4628 864
rect 4652 856 4660 864
rect 4412 816 4420 824
rect 4540 796 4548 804
rect 4556 776 4564 784
rect 4652 676 4660 684
rect 4684 676 4692 684
rect 4316 656 4324 664
rect 4380 616 4388 624
rect 4316 556 4324 564
rect 4348 556 4356 564
rect 4284 536 4292 544
rect 4268 496 4276 504
rect 4348 536 4356 544
rect 4396 516 4404 524
rect 4508 516 4516 524
rect 4332 496 4340 504
rect 4396 496 4404 504
rect 4444 496 4452 504
rect 4300 256 4308 264
rect 4012 156 4020 164
rect 4060 156 4068 164
rect 4108 156 4116 164
rect 4044 136 4052 144
rect 4044 116 4052 124
rect 4076 136 4084 144
rect 4172 136 4180 144
rect 4348 456 4356 464
rect 4364 316 4372 324
rect 4428 316 4436 324
rect 4508 476 4516 484
rect 4556 436 4564 444
rect 4460 316 4468 324
rect 4572 336 4580 344
rect 4428 296 4436 304
rect 4476 296 4484 304
rect 4364 256 4372 264
rect 4348 216 4356 224
rect 4300 196 4308 204
rect 4332 196 4340 204
rect 4316 156 4324 164
rect 4492 256 4500 264
rect 4524 256 4532 264
rect 4380 136 4388 144
rect 4428 136 4436 144
rect 4524 176 4532 184
rect 4684 656 4692 664
rect 4700 616 4708 624
rect 4668 456 4676 464
rect 5020 1318 5028 1324
rect 5244 1836 5252 1844
rect 5260 1836 5268 1844
rect 5228 1756 5236 1764
rect 5260 1796 5268 1804
rect 5324 1936 5332 1944
rect 5532 2156 5540 2164
rect 5804 2336 5812 2344
rect 5820 2336 5828 2344
rect 5676 2296 5684 2304
rect 5628 2276 5636 2284
rect 5644 2256 5652 2264
rect 5660 2256 5668 2264
rect 5612 2176 5620 2184
rect 5644 2156 5652 2164
rect 5548 2136 5556 2144
rect 5564 2116 5572 2124
rect 5692 2276 5700 2284
rect 5788 2276 5796 2284
rect 5724 2256 5732 2264
rect 5740 2256 5748 2264
rect 5692 2236 5700 2244
rect 5692 2156 5700 2164
rect 5788 2156 5796 2164
rect 5676 2116 5684 2124
rect 5724 2116 5732 2124
rect 5660 2096 5668 2104
rect 5916 2336 5924 2344
rect 5820 2296 5828 2304
rect 5836 2296 5844 2304
rect 5948 2396 5956 2404
rect 5932 2296 5940 2304
rect 5852 2276 5860 2284
rect 5900 2276 5908 2284
rect 5852 2156 5860 2164
rect 5916 2256 5924 2264
rect 5900 2236 5908 2244
rect 5884 2216 5892 2224
rect 5820 2116 5828 2124
rect 5900 2096 5908 2104
rect 5788 2076 5796 2084
rect 5868 2076 5876 2084
rect 5436 2036 5444 2044
rect 5580 2036 5588 2044
rect 5916 2036 5924 2044
rect 5756 1996 5764 2004
rect 5388 1916 5396 1924
rect 5468 1916 5476 1924
rect 5500 1916 5508 1924
rect 5660 1916 5668 1924
rect 5692 1916 5700 1924
rect 5340 1876 5348 1884
rect 5340 1816 5348 1824
rect 5372 1856 5380 1864
rect 5324 1796 5332 1804
rect 5356 1796 5364 1804
rect 5324 1756 5332 1764
rect 5420 1896 5428 1904
rect 5420 1876 5428 1884
rect 5468 1896 5476 1904
rect 5500 1896 5508 1904
rect 5548 1896 5556 1904
rect 5580 1896 5588 1904
rect 5692 1896 5700 1904
rect 5564 1876 5572 1884
rect 5644 1876 5652 1884
rect 5708 1876 5716 1884
rect 5516 1856 5524 1864
rect 5628 1856 5636 1864
rect 5724 1856 5732 1864
rect 5452 1816 5460 1824
rect 5468 1796 5476 1804
rect 5404 1776 5412 1784
rect 5308 1736 5316 1744
rect 5340 1736 5348 1744
rect 5436 1736 5444 1744
rect 5244 1716 5252 1724
rect 5260 1716 5268 1724
rect 5404 1676 5412 1684
rect 5260 1576 5268 1584
rect 5276 1556 5284 1564
rect 5228 1516 5236 1524
rect 5404 1556 5412 1564
rect 5228 1496 5236 1504
rect 5292 1496 5300 1504
rect 5340 1476 5348 1484
rect 5180 1456 5188 1464
rect 5340 1416 5348 1424
rect 5436 1396 5444 1404
rect 5388 1376 5396 1384
rect 5244 1356 5252 1364
rect 5276 1356 5284 1364
rect 5196 1336 5204 1344
rect 5452 1376 5460 1384
rect 5484 1436 5492 1444
rect 5500 1416 5508 1424
rect 5484 1376 5492 1384
rect 5484 1356 5492 1364
rect 5724 1836 5732 1844
rect 5532 1816 5540 1824
rect 5612 1796 5620 1804
rect 5660 1796 5668 1804
rect 5628 1756 5636 1764
rect 5708 1776 5716 1784
rect 5596 1716 5604 1724
rect 5836 1916 5844 1924
rect 5980 2356 5988 2364
rect 6108 2356 6116 2364
rect 5964 2256 5972 2264
rect 5948 1956 5956 1964
rect 5852 1896 5860 1904
rect 6268 2736 6276 2744
rect 6268 2696 6276 2704
rect 6748 3176 6756 3184
rect 6748 3156 6756 3164
rect 6508 3136 6516 3144
rect 6716 3136 6724 3144
rect 6460 3116 6468 3124
rect 6668 3116 6676 3124
rect 6588 3096 6596 3104
rect 6716 3096 6724 3104
rect 6396 3056 6404 3064
rect 6350 3006 6358 3014
rect 6364 3006 6372 3014
rect 6378 3006 6386 3014
rect 6348 2976 6356 2984
rect 6540 2976 6548 2984
rect 6476 2918 6484 2924
rect 6476 2916 6484 2918
rect 6636 3056 6644 3064
rect 6780 3096 6788 3104
rect 6812 3416 6820 3424
rect 6876 3496 6884 3504
rect 6924 3496 6932 3504
rect 6956 3496 6964 3504
rect 6876 3476 6884 3484
rect 6876 3416 6884 3424
rect 6860 3316 6868 3324
rect 7020 3736 7028 3744
rect 6988 3696 6996 3704
rect 7004 3556 7012 3564
rect 7084 3496 7092 3504
rect 6972 3436 6980 3444
rect 7052 3456 7060 3464
rect 7020 3416 7028 3424
rect 6908 3376 6916 3384
rect 6972 3376 6980 3384
rect 7068 3416 7076 3424
rect 7180 4136 7188 4144
rect 7228 4136 7236 4144
rect 7196 4116 7204 4124
rect 7244 4116 7252 4124
rect 7180 4096 7188 4104
rect 7164 4076 7172 4084
rect 7180 4016 7188 4024
rect 7132 3876 7140 3884
rect 7164 3876 7172 3884
rect 7388 4236 7396 4244
rect 7372 4216 7380 4224
rect 7372 4196 7380 4204
rect 7388 4156 7396 4164
rect 7276 4136 7284 4144
rect 7324 4136 7332 4144
rect 7372 4136 7380 4144
rect 7548 5456 7556 5464
rect 7484 5156 7492 5164
rect 7500 5116 7508 5124
rect 7564 5256 7572 5264
rect 7500 5076 7508 5084
rect 7484 5036 7492 5044
rect 7484 4696 7492 4704
rect 7484 4556 7492 4564
rect 7468 4536 7476 4544
rect 7452 4396 7460 4404
rect 7436 4356 7444 4364
rect 7436 4316 7444 4324
rect 7452 4296 7460 4304
rect 7516 4936 7524 4944
rect 7548 4918 7556 4924
rect 7548 4916 7556 4918
rect 7516 4756 7524 4764
rect 7532 4736 7540 4744
rect 7548 4696 7556 4704
rect 7564 4676 7572 4684
rect 7564 4616 7572 4624
rect 7596 5516 7604 5524
rect 7708 5636 7716 5644
rect 7756 5536 7764 5544
rect 8028 5718 8036 5724
rect 8028 5716 8036 5718
rect 8012 5636 8020 5644
rect 7836 5616 7844 5624
rect 7884 5556 7892 5564
rect 7948 5556 7956 5564
rect 7868 5536 7876 5544
rect 7916 5536 7924 5544
rect 7996 5536 8004 5544
rect 7852 5516 7860 5524
rect 7868 5496 7876 5504
rect 7900 5496 7908 5504
rect 7692 5476 7700 5484
rect 7820 5476 7828 5484
rect 7836 5456 7844 5464
rect 7628 5436 7636 5444
rect 7692 5436 7700 5444
rect 7708 5336 7716 5344
rect 7676 5236 7684 5244
rect 7676 5116 7684 5124
rect 7676 5096 7684 5104
rect 7756 5316 7764 5324
rect 7948 5456 7956 5464
rect 7948 5416 7956 5424
rect 7836 5336 7844 5344
rect 7868 5336 7876 5344
rect 7964 5356 7972 5364
rect 7900 5316 7908 5324
rect 7948 5316 7956 5324
rect 7740 5296 7748 5304
rect 7772 5296 7780 5304
rect 7788 5296 7796 5304
rect 7820 5296 7828 5304
rect 7772 5256 7780 5264
rect 7708 5136 7716 5144
rect 7740 5096 7748 5104
rect 7692 5076 7700 5084
rect 7740 5056 7748 5064
rect 7628 5016 7636 5024
rect 7724 5016 7732 5024
rect 7612 4996 7620 5004
rect 7772 4996 7780 5004
rect 7884 5296 7892 5304
rect 7804 5276 7812 5284
rect 7852 5276 7860 5284
rect 7820 5236 7828 5244
rect 7868 5236 7876 5244
rect 7804 5156 7812 5164
rect 7852 5156 7860 5164
rect 7852 5116 7860 5124
rect 7884 5136 7892 5144
rect 7916 5276 7924 5284
rect 7900 5116 7908 5124
rect 7932 5116 7940 5124
rect 7820 5076 7828 5084
rect 7852 5076 7860 5084
rect 7820 5056 7828 5064
rect 7820 5036 7828 5044
rect 7788 4956 7796 4964
rect 7676 4936 7684 4944
rect 7660 4916 7668 4924
rect 7724 4916 7732 4924
rect 7612 4876 7620 4884
rect 7644 4896 7652 4904
rect 7628 4836 7636 4844
rect 7596 4776 7604 4784
rect 7692 4896 7700 4904
rect 7724 4856 7732 4864
rect 7692 4836 7700 4844
rect 7708 4756 7716 4764
rect 7676 4736 7684 4744
rect 7692 4716 7700 4724
rect 7612 4676 7620 4684
rect 7628 4656 7636 4664
rect 7580 4596 7588 4604
rect 7564 4576 7572 4584
rect 7548 4556 7556 4564
rect 7660 4696 7668 4704
rect 7692 4696 7700 4704
rect 7676 4656 7684 4664
rect 7772 4916 7780 4924
rect 7772 4896 7780 4904
rect 7756 4736 7764 4744
rect 7836 4876 7844 4884
rect 7916 4976 7924 4984
rect 7948 4996 7956 5004
rect 7948 4976 7956 4984
rect 7932 4956 7940 4964
rect 7932 4936 7940 4944
rect 7868 4896 7876 4904
rect 7868 4796 7876 4804
rect 7852 4756 7860 4764
rect 7820 4716 7828 4724
rect 7804 4696 7812 4704
rect 7852 4696 7860 4704
rect 7820 4676 7828 4684
rect 7740 4656 7748 4664
rect 7788 4656 7796 4664
rect 7852 4656 7860 4664
rect 7724 4636 7732 4644
rect 7788 4636 7796 4644
rect 7692 4616 7700 4624
rect 7532 4536 7540 4544
rect 7644 4516 7652 4524
rect 7724 4556 7732 4564
rect 7772 4556 7780 4564
rect 7708 4536 7716 4544
rect 7484 4436 7492 4444
rect 7468 4276 7476 4284
rect 7436 4256 7444 4264
rect 7452 4256 7460 4264
rect 7436 4156 7444 4164
rect 7308 4116 7316 4124
rect 7324 4116 7332 4124
rect 7356 4116 7364 4124
rect 7308 3976 7316 3984
rect 7292 3936 7300 3944
rect 7404 4096 7412 4104
rect 7532 4416 7540 4424
rect 7500 4336 7508 4344
rect 7500 4236 7508 4244
rect 7468 4156 7476 4164
rect 7452 4076 7460 4084
rect 7468 4076 7476 4084
rect 7324 3896 7332 3904
rect 7356 3896 7364 3904
rect 7372 3896 7380 3904
rect 7468 3902 7476 3904
rect 7468 3896 7476 3902
rect 7580 4396 7588 4404
rect 7564 4356 7572 4364
rect 7628 4356 7636 4364
rect 7548 4296 7556 4304
rect 7596 4316 7604 4324
rect 7628 4296 7636 4304
rect 7580 4256 7588 4264
rect 7564 4196 7572 4204
rect 7692 4336 7700 4344
rect 7676 4256 7684 4264
rect 7644 4156 7652 4164
rect 7548 4116 7556 4124
rect 7612 4096 7620 4104
rect 7660 4096 7668 4104
rect 7612 4036 7620 4044
rect 7596 3976 7604 3984
rect 7612 3956 7620 3964
rect 7676 3916 7684 3924
rect 7564 3896 7572 3904
rect 7388 3876 7396 3884
rect 7532 3876 7540 3884
rect 7196 3856 7204 3864
rect 7260 3856 7268 3864
rect 7180 3756 7188 3764
rect 7148 3696 7156 3704
rect 7116 3676 7124 3684
rect 7164 3676 7172 3684
rect 7180 3556 7188 3564
rect 7148 3516 7156 3524
rect 7164 3476 7172 3484
rect 7100 3396 7108 3404
rect 7036 3376 7044 3384
rect 7068 3376 7076 3384
rect 7132 3376 7140 3384
rect 7372 3756 7380 3764
rect 7308 3736 7316 3744
rect 7212 3616 7220 3624
rect 7340 3696 7348 3704
rect 7324 3536 7332 3544
rect 7244 3516 7252 3524
rect 7084 3356 7092 3364
rect 7212 3356 7220 3364
rect 6892 3336 6900 3344
rect 6876 3176 6884 3184
rect 6860 3156 6868 3164
rect 6860 3116 6868 3124
rect 6844 3096 6852 3104
rect 6716 3036 6724 3044
rect 6684 3016 6692 3024
rect 6572 2956 6580 2964
rect 6636 2956 6644 2964
rect 6572 2936 6580 2944
rect 6620 2936 6628 2944
rect 6732 2996 6740 3004
rect 6588 2916 6596 2924
rect 6604 2916 6612 2924
rect 6700 2916 6708 2924
rect 6332 2876 6340 2884
rect 6508 2876 6516 2884
rect 6668 2876 6676 2884
rect 6300 2776 6308 2784
rect 6300 2696 6308 2704
rect 6284 2636 6292 2644
rect 6204 2616 6212 2624
rect 6236 2616 6244 2624
rect 6236 2596 6244 2604
rect 6204 2576 6212 2584
rect 6252 2556 6260 2564
rect 6236 2536 6244 2544
rect 6636 2696 6644 2704
rect 6796 3056 6804 3064
rect 6764 3016 6772 3024
rect 6876 3016 6884 3024
rect 6844 2996 6852 3004
rect 6844 2976 6852 2984
rect 7020 3316 7028 3324
rect 7260 3296 7268 3304
rect 7164 3276 7172 3284
rect 7292 3256 7300 3264
rect 7292 3236 7300 3244
rect 7084 3196 7092 3204
rect 7116 3196 7124 3204
rect 6972 3156 6980 3164
rect 6988 3156 6996 3164
rect 7036 3156 7044 3164
rect 6908 3116 6916 3124
rect 6940 3116 6948 3124
rect 7228 3136 7236 3144
rect 6972 3096 6980 3104
rect 7052 3096 7060 3104
rect 7004 3076 7012 3084
rect 6940 3056 6948 3064
rect 6988 3056 6996 3064
rect 7052 3056 7060 3064
rect 6924 2996 6932 3004
rect 6892 2956 6900 2964
rect 6908 2956 6916 2964
rect 6764 2918 6772 2924
rect 6764 2916 6772 2918
rect 6860 2916 6868 2924
rect 6780 2696 6788 2704
rect 6988 3016 6996 3024
rect 7036 3016 7044 3024
rect 6972 2996 6980 3004
rect 6956 2976 6964 2984
rect 6940 2936 6948 2944
rect 6924 2916 6932 2924
rect 6940 2896 6948 2904
rect 7132 3096 7140 3104
rect 7180 3096 7188 3104
rect 7260 3096 7268 3104
rect 7292 3096 7300 3104
rect 7180 3076 7188 3084
rect 7228 3076 7236 3084
rect 7148 3036 7156 3044
rect 7132 3016 7140 3024
rect 6956 2776 6964 2784
rect 6988 2776 6996 2784
rect 7340 3056 7348 3064
rect 7372 2956 7380 2964
rect 7404 3856 7412 3864
rect 7436 3736 7444 3744
rect 7452 3736 7460 3744
rect 7468 3716 7476 3724
rect 7532 3756 7540 3764
rect 7548 3736 7556 3744
rect 7484 3696 7492 3704
rect 7500 3696 7508 3704
rect 7420 3676 7428 3684
rect 7596 3736 7604 3744
rect 7660 3756 7668 3764
rect 7708 4156 7716 4164
rect 7708 4136 7716 4144
rect 7852 4536 7860 4544
rect 7836 4516 7844 4524
rect 7756 4336 7764 4344
rect 7772 4336 7780 4344
rect 7804 4336 7812 4344
rect 7740 4316 7748 4324
rect 7772 4296 7780 4304
rect 7788 4216 7796 4224
rect 7756 4176 7764 4184
rect 7740 4076 7748 4084
rect 7788 4076 7796 4084
rect 7820 4316 7828 4324
rect 7836 4296 7844 4304
rect 7820 4276 7828 4284
rect 7804 4056 7812 4064
rect 7772 4036 7780 4044
rect 7804 4036 7812 4044
rect 7996 5416 8004 5424
rect 8076 5516 8084 5524
rect 8076 5496 8084 5504
rect 8124 5496 8132 5504
rect 8108 5476 8116 5484
rect 8044 5436 8052 5444
rect 8028 5376 8036 5384
rect 8076 5376 8084 5384
rect 8140 5356 8148 5364
rect 7980 5336 7988 5344
rect 8028 5336 8036 5344
rect 7996 5316 8004 5324
rect 8044 5316 8052 5324
rect 8140 5316 8148 5324
rect 8028 5296 8036 5304
rect 7980 5276 7988 5284
rect 8012 5276 8020 5284
rect 8060 5116 8068 5124
rect 8076 5116 8084 5124
rect 8044 5096 8052 5104
rect 8028 5076 8036 5084
rect 8012 5056 8020 5064
rect 7996 5036 8004 5044
rect 7980 5016 7988 5024
rect 7996 4956 8004 4964
rect 7964 4876 7972 4884
rect 7900 4856 7908 4864
rect 7884 4736 7892 4744
rect 7884 4676 7892 4684
rect 7964 4796 7972 4804
rect 7948 4696 7956 4704
rect 7916 4676 7924 4684
rect 7916 4656 7924 4664
rect 8044 4876 8052 4884
rect 8092 5096 8100 5104
rect 8092 4936 8100 4944
rect 8124 4916 8132 4924
rect 8124 4876 8132 4884
rect 8108 4856 8116 4864
rect 8092 4756 8100 4764
rect 8060 4736 8068 4744
rect 7996 4716 8004 4724
rect 8060 4716 8068 4724
rect 8012 4696 8020 4704
rect 7900 4616 7908 4624
rect 7916 4536 7924 4544
rect 7900 4356 7908 4364
rect 8028 4656 8036 4664
rect 8076 4636 8084 4644
rect 8044 4616 8052 4624
rect 7996 4596 8004 4604
rect 8028 4596 8036 4604
rect 8012 4536 8020 4544
rect 7980 4516 7988 4524
rect 7932 4476 7940 4484
rect 7836 4156 7844 4164
rect 7836 4036 7844 4044
rect 7820 4016 7828 4024
rect 7740 3956 7748 3964
rect 7788 3956 7796 3964
rect 7708 3916 7716 3924
rect 7708 3896 7716 3904
rect 7724 3856 7732 3864
rect 7644 3736 7652 3744
rect 7644 3716 7652 3724
rect 7612 3696 7620 3704
rect 7628 3696 7636 3704
rect 7580 3656 7588 3664
rect 7564 3516 7572 3524
rect 7596 3516 7604 3524
rect 7724 3516 7732 3524
rect 7484 3496 7492 3504
rect 7516 3496 7524 3504
rect 7436 3456 7444 3464
rect 7644 3476 7652 3484
rect 7660 3456 7668 3464
rect 7692 3456 7700 3464
rect 7500 3336 7508 3344
rect 7516 3336 7524 3344
rect 7500 3316 7508 3324
rect 7420 3276 7428 3284
rect 7532 3316 7540 3324
rect 7548 3316 7556 3324
rect 7612 3316 7620 3324
rect 7676 3396 7684 3404
rect 7708 3396 7716 3404
rect 7676 3336 7684 3344
rect 7516 3296 7524 3304
rect 7596 3296 7604 3304
rect 7612 3296 7620 3304
rect 7532 3276 7540 3284
rect 7484 3176 7492 3184
rect 7452 3156 7460 3164
rect 7484 3156 7492 3164
rect 7628 3256 7636 3264
rect 7500 3116 7508 3124
rect 7532 3116 7540 3124
rect 7612 3116 7620 3124
rect 7452 3056 7460 3064
rect 7580 3096 7588 3104
rect 7628 3096 7636 3104
rect 7660 3276 7668 3284
rect 7660 3096 7668 3104
rect 7596 3076 7604 3084
rect 7644 3076 7652 3084
rect 7692 3296 7700 3304
rect 7724 3356 7732 3364
rect 7756 3856 7764 3864
rect 7756 3716 7764 3724
rect 7788 3716 7796 3724
rect 7788 3656 7796 3664
rect 7772 3516 7780 3524
rect 7836 3736 7844 3744
rect 7820 3716 7828 3724
rect 7900 4116 7908 4124
rect 7868 4056 7876 4064
rect 7900 4056 7908 4064
rect 7884 3996 7892 4004
rect 7884 3976 7892 3984
rect 7868 3896 7876 3904
rect 7868 3756 7876 3764
rect 7948 4396 7956 4404
rect 8060 4516 8068 4524
rect 8060 4396 8068 4404
rect 7964 4256 7972 4264
rect 8028 4196 8036 4204
rect 7948 4176 7956 4184
rect 8012 4136 8020 4144
rect 7964 4076 7972 4084
rect 7964 4056 7972 4064
rect 7932 3936 7940 3944
rect 7948 3916 7956 3924
rect 7948 3896 7956 3904
rect 7948 3856 7956 3864
rect 8012 4076 8020 4084
rect 7996 3976 8004 3984
rect 7980 3956 7988 3964
rect 7996 3956 8004 3964
rect 7980 3876 7988 3884
rect 8012 3836 8020 3844
rect 7916 3716 7924 3724
rect 7900 3676 7908 3684
rect 7820 3656 7828 3664
rect 7852 3656 7860 3664
rect 7772 3496 7780 3504
rect 7804 3496 7812 3504
rect 7756 3376 7764 3384
rect 7740 3316 7748 3324
rect 7788 3396 7796 3404
rect 7756 3296 7764 3304
rect 7772 3296 7780 3304
rect 7692 3276 7700 3284
rect 7900 3516 7908 3524
rect 7980 3476 7988 3484
rect 7980 3436 7988 3444
rect 7836 3356 7844 3364
rect 7948 3356 7956 3364
rect 7852 3336 7860 3344
rect 7884 3316 7892 3324
rect 7996 3316 8004 3324
rect 7964 3296 7972 3304
rect 7820 3276 7828 3284
rect 7852 3276 7860 3284
rect 7804 3256 7812 3264
rect 7724 3216 7732 3224
rect 7788 3216 7796 3224
rect 7788 3136 7796 3144
rect 7804 3116 7812 3124
rect 7740 3096 7748 3104
rect 7836 3156 7844 3164
rect 7548 3056 7556 3064
rect 7564 3056 7572 3064
rect 7628 3036 7636 3044
rect 7420 2996 7428 3004
rect 7516 2996 7524 3004
rect 7676 2996 7684 3004
rect 7724 2996 7732 3004
rect 7708 2976 7716 2984
rect 7436 2956 7444 2964
rect 7500 2956 7508 2964
rect 7660 2956 7668 2964
rect 7036 2936 7044 2944
rect 7356 2936 7364 2944
rect 7036 2916 7044 2924
rect 7068 2916 7076 2924
rect 7084 2916 7092 2924
rect 7132 2916 7140 2924
rect 7052 2696 7060 2704
rect 7148 2816 7156 2824
rect 7180 2796 7188 2804
rect 7324 2796 7332 2804
rect 7148 2716 7156 2724
rect 6508 2676 6516 2684
rect 6652 2676 6660 2684
rect 6716 2676 6724 2684
rect 6350 2606 6358 2614
rect 6364 2606 6372 2614
rect 6378 2606 6386 2614
rect 6428 2636 6436 2644
rect 6412 2576 6420 2584
rect 6348 2556 6356 2564
rect 6444 2556 6452 2564
rect 6748 2616 6756 2624
rect 6764 2596 6772 2604
rect 6524 2536 6532 2544
rect 6588 2536 6596 2544
rect 6780 2536 6788 2544
rect 6252 2516 6260 2524
rect 6364 2516 6372 2524
rect 6204 2496 6212 2504
rect 6268 2496 6276 2504
rect 6300 2476 6308 2484
rect 6220 2456 6228 2464
rect 6284 2356 6292 2364
rect 6060 2316 6068 2324
rect 6124 2336 6132 2344
rect 6188 2336 6196 2344
rect 6540 2476 6548 2484
rect 6204 2316 6212 2324
rect 6316 2316 6324 2324
rect 6428 2316 6436 2324
rect 6620 2516 6628 2524
rect 6684 2516 6692 2524
rect 6812 2518 6820 2524
rect 6812 2516 6820 2518
rect 6604 2476 6612 2484
rect 6668 2476 6676 2484
rect 6300 2296 6308 2304
rect 6076 2276 6084 2284
rect 6108 2276 6116 2284
rect 6012 2216 6020 2224
rect 6028 2156 6036 2164
rect 6044 2156 6052 2164
rect 6076 2156 6084 2164
rect 6172 2276 6180 2284
rect 6204 2276 6212 2284
rect 6460 2276 6468 2284
rect 6156 2236 6164 2244
rect 6172 2176 6180 2184
rect 6252 2256 6260 2264
rect 6332 2256 6340 2264
rect 6236 2156 6244 2164
rect 6076 2136 6084 2144
rect 6220 2136 6228 2144
rect 6108 2076 6116 2084
rect 6412 2236 6420 2244
rect 6350 2206 6358 2214
rect 6364 2206 6372 2214
rect 6378 2206 6386 2214
rect 6332 2176 6340 2184
rect 6284 2156 6292 2164
rect 6540 2236 6548 2244
rect 6524 2196 6532 2204
rect 6860 2376 6868 2384
rect 6668 2356 6676 2364
rect 6764 2356 6772 2364
rect 6748 2296 6756 2304
rect 6652 2236 6660 2244
rect 6652 2216 6660 2224
rect 6476 2156 6484 2164
rect 6540 2156 6548 2164
rect 6572 2156 6580 2164
rect 6364 2136 6372 2144
rect 6444 2116 6452 2124
rect 6316 2096 6324 2104
rect 6444 2096 6452 2104
rect 6524 2096 6532 2104
rect 6476 2056 6484 2064
rect 6252 2016 6260 2024
rect 6076 1956 6084 1964
rect 6028 1896 6036 1904
rect 5980 1836 5988 1844
rect 5948 1776 5956 1784
rect 5756 1756 5764 1764
rect 5884 1756 5892 1764
rect 5932 1756 5940 1764
rect 6012 1756 6020 1764
rect 5788 1736 5796 1744
rect 5820 1718 5828 1724
rect 5820 1716 5828 1718
rect 6172 1896 6180 1904
rect 6092 1836 6100 1844
rect 6124 1836 6132 1844
rect 5692 1576 5700 1584
rect 5708 1556 5716 1564
rect 5692 1536 5700 1544
rect 5548 1516 5556 1524
rect 5980 1536 5988 1544
rect 5628 1496 5636 1504
rect 5596 1476 5604 1484
rect 5532 1396 5540 1404
rect 5276 1336 5284 1344
rect 5308 1336 5316 1344
rect 5468 1336 5476 1344
rect 5516 1336 5524 1344
rect 5020 1316 5028 1318
rect 4876 1276 4884 1284
rect 4940 1276 4948 1284
rect 4860 1256 4868 1264
rect 4814 1206 4822 1214
rect 4828 1206 4836 1214
rect 4842 1206 4850 1214
rect 4796 1156 4804 1164
rect 4796 1076 4804 1084
rect 4780 956 4788 964
rect 4796 956 4804 964
rect 4780 896 4788 904
rect 4988 1256 4996 1264
rect 4908 1096 4916 1104
rect 4924 1096 4932 1104
rect 4892 1080 4900 1084
rect 4892 1076 4900 1080
rect 4908 1056 4916 1064
rect 4908 976 4916 984
rect 4812 936 4820 944
rect 4796 856 4804 864
rect 5068 1196 5076 1204
rect 4956 1116 4964 1124
rect 4988 1116 4996 1124
rect 5052 1116 5060 1124
rect 5004 1096 5012 1104
rect 4988 1056 4996 1064
rect 4940 1016 4948 1024
rect 5068 1076 5076 1084
rect 5020 1056 5028 1064
rect 5020 1016 5028 1024
rect 5004 996 5012 1004
rect 5116 1076 5124 1084
rect 5084 1056 5092 1064
rect 5100 1056 5108 1064
rect 5068 976 5076 984
rect 5052 956 5060 964
rect 5100 1016 5108 1024
rect 4972 936 4980 944
rect 4972 916 4980 924
rect 5164 1316 5172 1324
rect 5196 1316 5204 1324
rect 5244 1316 5252 1324
rect 5276 1316 5284 1324
rect 5148 1296 5156 1304
rect 5212 1276 5220 1284
rect 5148 1216 5156 1224
rect 5436 1256 5444 1264
rect 5324 1236 5332 1244
rect 5308 1216 5316 1224
rect 5164 1176 5172 1184
rect 5164 1116 5172 1124
rect 5244 1116 5252 1124
rect 5148 1076 5156 1084
rect 5180 1096 5188 1104
rect 5212 1096 5220 1104
rect 5244 1096 5252 1104
rect 5260 1096 5268 1104
rect 5180 1036 5188 1044
rect 5228 1016 5236 1024
rect 5276 1076 5284 1084
rect 5292 1076 5300 1084
rect 5260 996 5268 1004
rect 5212 976 5220 984
rect 5292 956 5300 964
rect 4924 896 4932 904
rect 4956 896 4964 904
rect 5132 896 5140 904
rect 4892 856 4900 864
rect 4844 836 4852 844
rect 4860 836 4868 844
rect 4814 806 4822 814
rect 4828 806 4836 814
rect 4842 806 4850 814
rect 4780 696 4788 704
rect 4844 702 4852 704
rect 4844 696 4852 702
rect 4876 656 4884 664
rect 4908 616 4916 624
rect 5212 876 5220 884
rect 4988 836 4996 844
rect 5132 756 5140 764
rect 5196 756 5204 764
rect 5132 736 5140 744
rect 5068 716 5076 724
rect 5100 716 5108 724
rect 5180 716 5188 724
rect 5068 696 5076 704
rect 4988 676 4996 684
rect 4972 636 4980 644
rect 5004 636 5012 644
rect 5084 616 5092 624
rect 5228 736 5236 744
rect 5148 676 5156 684
rect 5148 616 5156 624
rect 4780 556 4788 564
rect 4924 556 4932 564
rect 4956 556 4964 564
rect 4892 536 4900 544
rect 4972 536 4980 544
rect 5004 536 5012 544
rect 5052 536 5060 544
rect 4764 516 4772 524
rect 4796 516 4804 524
rect 4814 406 4822 414
rect 4828 406 4836 414
rect 4842 406 4850 414
rect 4940 356 4948 364
rect 4940 336 4948 344
rect 4588 316 4596 324
rect 4620 316 4628 324
rect 4636 316 4644 324
rect 4604 296 4612 304
rect 4572 216 4580 224
rect 4508 156 4516 164
rect 4540 156 4548 164
rect 4588 156 4596 164
rect 4556 136 4564 144
rect 4572 136 4580 144
rect 4636 296 4644 304
rect 4652 296 4660 304
rect 4700 316 4708 324
rect 4652 256 4660 264
rect 4684 256 4692 264
rect 4620 216 4628 224
rect 4732 296 4740 304
rect 4684 176 4692 184
rect 4716 176 4724 184
rect 4636 136 4644 144
rect 4796 236 4804 244
rect 4812 176 4820 184
rect 4732 156 4740 164
rect 4764 136 4772 144
rect 4860 236 4868 244
rect 4844 156 4852 164
rect 4876 216 4884 224
rect 4892 216 4900 224
rect 4988 516 4996 524
rect 5132 596 5140 604
rect 5388 1196 5396 1204
rect 5340 1156 5348 1164
rect 5372 1116 5380 1124
rect 5404 1156 5412 1164
rect 5340 1096 5348 1104
rect 5356 1076 5364 1084
rect 5420 1076 5428 1084
rect 5436 1036 5444 1044
rect 5388 936 5396 944
rect 5580 1396 5588 1404
rect 5628 1396 5636 1404
rect 5580 1376 5588 1384
rect 5548 1336 5556 1344
rect 5756 1496 5764 1504
rect 5772 1496 5780 1504
rect 5804 1496 5812 1504
rect 5820 1496 5828 1504
rect 5820 1476 5828 1484
rect 5884 1476 5892 1484
rect 5932 1476 5940 1484
rect 5772 1416 5780 1424
rect 5756 1376 5764 1384
rect 5788 1376 5796 1384
rect 5660 1356 5668 1364
rect 5740 1356 5748 1364
rect 5724 1316 5732 1324
rect 5772 1316 5780 1324
rect 5644 1296 5652 1304
rect 5692 1296 5700 1304
rect 5676 1256 5684 1264
rect 5612 1236 5620 1244
rect 5708 1236 5716 1244
rect 5756 1236 5764 1244
rect 5516 1156 5524 1164
rect 5628 1136 5636 1144
rect 5532 1076 5540 1084
rect 5708 1116 5716 1124
rect 5676 1096 5684 1104
rect 5708 1096 5716 1104
rect 5596 1056 5604 1064
rect 5484 956 5492 964
rect 5628 1036 5636 1044
rect 5644 996 5652 1004
rect 5532 936 5540 944
rect 5564 936 5572 944
rect 5356 918 5364 924
rect 5356 916 5364 918
rect 5468 916 5476 924
rect 5308 876 5316 884
rect 5420 876 5428 884
rect 5852 1436 5860 1444
rect 5900 1396 5908 1404
rect 5964 1396 5972 1404
rect 6140 1776 6148 1784
rect 6268 1936 6276 1944
rect 6284 1916 6292 1924
rect 6412 1916 6420 1924
rect 6732 2236 6740 2244
rect 6956 2636 6964 2644
rect 6940 2616 6948 2624
rect 6972 2376 6980 2384
rect 6924 2356 6932 2364
rect 7004 2356 7012 2364
rect 6908 2336 6916 2344
rect 6796 2316 6804 2324
rect 6876 2316 6884 2324
rect 6892 2296 6900 2304
rect 6988 2316 6996 2324
rect 6940 2296 6948 2304
rect 6988 2296 6996 2304
rect 6860 2276 6868 2284
rect 6764 2236 6772 2244
rect 6812 2236 6820 2244
rect 6700 2196 6708 2204
rect 6684 2176 6692 2184
rect 6700 2176 6708 2184
rect 6732 2156 6740 2164
rect 6748 2156 6756 2164
rect 6700 2136 6708 2144
rect 6716 2096 6724 2104
rect 6716 2076 6724 2084
rect 6668 2056 6676 2064
rect 6636 2036 6644 2044
rect 6668 2036 6676 2044
rect 6588 1996 6596 2004
rect 6556 1936 6564 1944
rect 6332 1896 6340 1904
rect 6412 1896 6420 1904
rect 6492 1896 6500 1904
rect 6524 1896 6532 1904
rect 6252 1836 6260 1844
rect 6444 1856 6452 1864
rect 6350 1806 6358 1814
rect 6364 1806 6372 1814
rect 6378 1806 6386 1814
rect 6524 1876 6532 1884
rect 6572 1876 6580 1884
rect 6588 1856 6596 1864
rect 6604 1856 6612 1864
rect 6460 1836 6468 1844
rect 6444 1776 6452 1784
rect 6396 1756 6404 1764
rect 6476 1756 6484 1764
rect 6364 1736 6372 1744
rect 6172 1676 6180 1684
rect 6156 1596 6164 1604
rect 6108 1556 6116 1564
rect 6124 1536 6132 1544
rect 5868 1356 5876 1364
rect 5884 1356 5892 1364
rect 6044 1356 6052 1364
rect 5868 1256 5876 1264
rect 5836 1236 5844 1244
rect 5820 1196 5828 1204
rect 5788 1116 5796 1124
rect 5948 1236 5956 1244
rect 5900 1156 5908 1164
rect 5868 1116 5876 1124
rect 5916 1116 5924 1124
rect 5932 1096 5940 1104
rect 5980 1136 5988 1144
rect 5916 1076 5924 1084
rect 5772 1056 5780 1064
rect 5724 996 5732 1004
rect 5852 996 5860 1004
rect 6332 1656 6340 1664
rect 6268 1616 6276 1624
rect 6252 1536 6260 1544
rect 6220 1496 6228 1504
rect 6300 1496 6308 1504
rect 6524 1776 6532 1784
rect 6572 1776 6580 1784
rect 6540 1756 6548 1764
rect 6636 1836 6644 1844
rect 6588 1756 6596 1764
rect 6620 1756 6628 1764
rect 6492 1736 6500 1744
rect 6508 1736 6516 1744
rect 6604 1736 6612 1744
rect 6444 1716 6452 1724
rect 6524 1716 6532 1724
rect 6428 1656 6436 1664
rect 6476 1696 6484 1704
rect 6492 1696 6500 1704
rect 6588 1696 6596 1704
rect 6636 1676 6644 1684
rect 6716 1876 6724 1884
rect 6780 2216 6788 2224
rect 6796 2156 6804 2164
rect 6780 2136 6788 2144
rect 6844 2176 6852 2184
rect 6860 2136 6868 2144
rect 6924 2216 6932 2224
rect 6892 2116 6900 2124
rect 6908 2116 6916 2124
rect 6748 2096 6756 2104
rect 6764 2076 6772 2084
rect 6844 2096 6852 2104
rect 6908 2096 6916 2104
rect 6876 2076 6884 2084
rect 6812 2056 6820 2064
rect 6780 1916 6788 1924
rect 6764 1896 6772 1904
rect 6876 1996 6884 2004
rect 6844 1896 6852 1904
rect 6844 1876 6852 1884
rect 6796 1856 6804 1864
rect 6732 1836 6740 1844
rect 6812 1796 6820 1804
rect 6684 1776 6692 1784
rect 6700 1776 6708 1784
rect 6668 1736 6676 1744
rect 6588 1656 6596 1664
rect 6652 1656 6660 1664
rect 6460 1596 6468 1604
rect 6476 1596 6484 1604
rect 6428 1576 6436 1584
rect 6396 1556 6404 1564
rect 6412 1496 6420 1504
rect 6284 1476 6292 1484
rect 6124 1456 6132 1464
rect 6188 1456 6196 1464
rect 6204 1456 6212 1464
rect 6236 1456 6244 1464
rect 6108 1396 6116 1404
rect 6124 1356 6132 1364
rect 6156 1336 6164 1344
rect 6350 1406 6358 1414
rect 6364 1406 6372 1414
rect 6378 1406 6386 1414
rect 6284 1376 6292 1384
rect 6188 1316 6196 1324
rect 6220 1318 6228 1324
rect 6220 1316 6228 1318
rect 6156 1296 6164 1304
rect 6060 1216 6068 1224
rect 6028 1076 6036 1084
rect 5708 956 5716 964
rect 5996 956 6004 964
rect 5692 936 5700 944
rect 5676 916 5684 924
rect 5660 896 5668 904
rect 5516 816 5524 824
rect 5612 816 5620 824
rect 5564 736 5572 744
rect 5532 716 5540 724
rect 5340 696 5348 704
rect 5580 696 5588 704
rect 5292 676 5300 684
rect 5484 676 5492 684
rect 5388 656 5396 664
rect 5436 656 5444 664
rect 5180 556 5188 564
rect 5100 516 5108 524
rect 5036 496 5044 504
rect 5084 476 5092 484
rect 5100 456 5108 464
rect 5020 356 5028 364
rect 5100 356 5108 364
rect 5068 336 5076 344
rect 4988 316 4996 324
rect 4924 176 4932 184
rect 4924 156 4932 164
rect 5068 296 5076 304
rect 5084 256 5092 264
rect 5116 336 5124 344
rect 5132 336 5140 344
rect 5196 536 5204 544
rect 5468 636 5476 644
rect 5452 556 5460 564
rect 5484 536 5492 544
rect 5564 596 5572 604
rect 5564 556 5572 564
rect 5340 516 5348 524
rect 5532 516 5540 524
rect 5260 496 5268 504
rect 5196 376 5204 384
rect 5132 176 5140 184
rect 5164 296 5172 304
rect 5244 476 5252 484
rect 5228 336 5236 344
rect 5228 296 5236 304
rect 5196 256 5204 264
rect 5212 256 5220 264
rect 5148 156 5156 164
rect 5020 136 5028 144
rect 5164 136 5172 144
rect 5228 216 5236 224
rect 5212 156 5220 164
rect 5212 136 5220 144
rect 5308 376 5316 384
rect 5276 296 5284 304
rect 5628 536 5636 544
rect 5420 416 5428 424
rect 5452 396 5460 404
rect 5388 356 5396 364
rect 5532 356 5540 364
rect 5484 296 5492 304
rect 5292 256 5300 264
rect 5340 256 5348 264
rect 5260 176 5268 184
rect 5308 156 5316 164
rect 5484 216 5492 224
rect 5372 176 5380 184
rect 5468 176 5476 184
rect 5596 496 5604 504
rect 5612 456 5620 464
rect 5772 936 5780 944
rect 6108 1176 6116 1184
rect 6076 1116 6084 1124
rect 6204 1196 6212 1204
rect 6172 1096 6180 1104
rect 6188 1096 6196 1104
rect 6220 1176 6228 1184
rect 6236 1116 6244 1124
rect 6268 1116 6276 1124
rect 6268 1096 6276 1104
rect 6092 1056 6100 1064
rect 6204 1016 6212 1024
rect 6268 976 6276 984
rect 6060 936 6068 944
rect 6124 936 6132 944
rect 6540 1536 6548 1544
rect 6508 1496 6516 1504
rect 6572 1496 6580 1504
rect 6540 1476 6548 1484
rect 6572 1416 6580 1424
rect 6460 1376 6468 1384
rect 6556 1376 6564 1384
rect 6444 1356 6452 1364
rect 6460 1356 6468 1364
rect 6620 1616 6628 1624
rect 6652 1476 6660 1484
rect 6620 1456 6628 1464
rect 6732 1756 6740 1764
rect 6828 1756 6836 1764
rect 6700 1676 6708 1684
rect 6748 1716 6756 1724
rect 7036 2336 7044 2344
rect 7116 2556 7124 2564
rect 7404 2916 7412 2924
rect 7484 2916 7492 2924
rect 7388 2776 7396 2784
rect 7420 2756 7428 2764
rect 7356 2736 7364 2744
rect 7404 2716 7412 2724
rect 7468 2896 7476 2904
rect 7788 3036 7796 3044
rect 7836 2976 7844 2984
rect 7596 2936 7604 2944
rect 7484 2776 7492 2784
rect 7516 2716 7524 2724
rect 7628 2896 7636 2904
rect 7564 2716 7572 2724
rect 7212 2696 7220 2704
rect 7260 2696 7268 2704
rect 7452 2696 7460 2704
rect 7596 2696 7604 2704
rect 7228 2536 7236 2544
rect 7084 2518 7092 2524
rect 7084 2516 7092 2518
rect 7212 2516 7220 2524
rect 7180 2496 7188 2504
rect 7244 2496 7252 2504
rect 7340 2676 7348 2684
rect 7372 2656 7380 2664
rect 7308 2636 7316 2644
rect 7276 2576 7284 2584
rect 7356 2556 7364 2564
rect 7340 2518 7348 2524
rect 7340 2516 7348 2518
rect 7100 2336 7108 2344
rect 7228 2336 7236 2344
rect 7068 2156 7076 2164
rect 7004 2136 7012 2144
rect 7052 2116 7060 2124
rect 7276 2456 7284 2464
rect 7116 2316 7124 2324
rect 7116 2176 7124 2184
rect 7132 2136 7140 2144
rect 7148 2136 7156 2144
rect 6956 2096 6964 2104
rect 7036 2096 7044 2104
rect 6924 2016 6932 2024
rect 6924 1916 6932 1924
rect 7020 1916 7028 1924
rect 6892 1896 6900 1904
rect 6988 1902 6996 1904
rect 6988 1896 6996 1902
rect 7020 1876 7028 1884
rect 6876 1856 6884 1864
rect 6988 1856 6996 1864
rect 6892 1796 6900 1804
rect 6892 1776 6900 1784
rect 6972 1716 6980 1724
rect 6860 1696 6868 1704
rect 6972 1696 6980 1704
rect 6876 1676 6884 1684
rect 6780 1656 6788 1664
rect 6876 1636 6884 1644
rect 7148 2076 7156 2084
rect 7068 1996 7076 2004
rect 7212 2176 7220 2184
rect 7180 2156 7188 2164
rect 7244 2296 7252 2304
rect 7356 2436 7364 2444
rect 7340 2356 7348 2364
rect 7420 2676 7428 2684
rect 7452 2656 7460 2664
rect 7388 2636 7396 2644
rect 7740 2916 7748 2924
rect 7788 2916 7796 2924
rect 7484 2676 7492 2684
rect 7580 2676 7588 2684
rect 7676 2676 7684 2684
rect 7468 2576 7476 2584
rect 7532 2656 7540 2664
rect 7580 2656 7588 2664
rect 7516 2596 7524 2604
rect 7564 2596 7572 2604
rect 7500 2516 7508 2524
rect 7644 2596 7652 2604
rect 7676 2636 7684 2644
rect 7836 2896 7844 2904
rect 7836 2856 7844 2864
rect 7804 2776 7812 2784
rect 7804 2696 7812 2704
rect 8044 4176 8052 4184
rect 8044 4156 8052 4164
rect 8124 4616 8132 4624
rect 8092 4436 8100 4444
rect 8076 4196 8084 4204
rect 8076 4136 8084 4144
rect 8044 4036 8052 4044
rect 8108 4116 8116 4124
rect 8092 4096 8100 4104
rect 8092 4016 8100 4024
rect 8092 3996 8100 4004
rect 8108 3956 8116 3964
rect 8060 3916 8068 3924
rect 8044 3896 8052 3904
rect 8092 3896 8100 3904
rect 8060 3856 8068 3864
rect 8108 3776 8116 3784
rect 8108 3736 8116 3744
rect 8044 3716 8052 3724
rect 8092 3716 8100 3724
rect 8108 3716 8116 3724
rect 8076 3556 8084 3564
rect 8044 3496 8052 3504
rect 7948 3176 7956 3184
rect 8012 3176 8020 3184
rect 8028 3156 8036 3164
rect 7932 3136 7940 3144
rect 7868 3116 7876 3124
rect 7900 3116 7908 3124
rect 8028 3116 8036 3124
rect 7868 3076 7876 3084
rect 7884 2876 7892 2884
rect 8012 3096 8020 3104
rect 7916 3056 7924 3064
rect 7932 2956 7940 2964
rect 7932 2896 7940 2904
rect 7900 2856 7908 2864
rect 7932 2856 7940 2864
rect 7868 2736 7876 2744
rect 7900 2736 7908 2744
rect 7996 2916 8004 2924
rect 7964 2736 7972 2744
rect 8012 2756 8020 2764
rect 7916 2696 7924 2704
rect 7948 2696 7956 2704
rect 7852 2676 7860 2684
rect 7836 2656 7844 2664
rect 7948 2676 7956 2684
rect 7868 2656 7876 2664
rect 7964 2656 7972 2664
rect 7852 2636 7860 2644
rect 7788 2616 7796 2624
rect 7660 2556 7668 2564
rect 7740 2556 7748 2564
rect 7548 2536 7556 2544
rect 7580 2516 7588 2524
rect 7484 2436 7492 2444
rect 7420 2376 7428 2384
rect 7404 2316 7412 2324
rect 7244 2116 7252 2124
rect 7148 1876 7156 1884
rect 7196 1876 7204 1884
rect 7116 1836 7124 1844
rect 7292 2216 7300 2224
rect 7276 2196 7284 2204
rect 7308 2196 7316 2204
rect 7276 2176 7284 2184
rect 7292 2176 7300 2184
rect 7516 2376 7524 2384
rect 7516 2336 7524 2344
rect 7500 2296 7508 2304
rect 7468 2276 7476 2284
rect 7628 2516 7636 2524
rect 7612 2436 7620 2444
rect 7564 2316 7572 2324
rect 7580 2316 7588 2324
rect 7596 2296 7604 2304
rect 7676 2516 7684 2524
rect 7708 2516 7716 2524
rect 7740 2516 7748 2524
rect 7740 2356 7748 2364
rect 7740 2336 7748 2344
rect 7804 2516 7812 2524
rect 7836 2516 7844 2524
rect 7788 2476 7796 2484
rect 7772 2356 7780 2364
rect 7804 2336 7812 2344
rect 7756 2316 7764 2324
rect 7788 2316 7796 2324
rect 7660 2296 7668 2304
rect 7724 2296 7732 2304
rect 7788 2296 7796 2304
rect 7820 2296 7828 2304
rect 7452 2256 7460 2264
rect 7516 2256 7524 2264
rect 7612 2256 7620 2264
rect 7388 2176 7396 2184
rect 7372 2156 7380 2164
rect 7468 2156 7476 2164
rect 7324 2136 7332 2144
rect 7420 2136 7428 2144
rect 7228 2096 7236 2104
rect 7356 2096 7364 2104
rect 7276 1976 7284 1984
rect 7324 1976 7332 1984
rect 7308 1956 7316 1964
rect 7324 1916 7332 1924
rect 7276 1896 7284 1904
rect 7420 1896 7428 1904
rect 7260 1796 7268 1804
rect 7212 1776 7220 1784
rect 7116 1756 7124 1764
rect 7180 1756 7188 1764
rect 7324 1876 7332 1884
rect 7084 1716 7092 1724
rect 7452 1916 7460 1924
rect 7580 2176 7588 2184
rect 7500 2136 7508 2144
rect 7548 2136 7556 2144
rect 7740 2136 7748 2144
rect 7852 2296 7860 2304
rect 7852 2276 7860 2284
rect 7836 2256 7844 2264
rect 7500 2116 7508 2124
rect 7708 2118 7716 2124
rect 7708 2116 7716 2118
rect 7788 2116 7796 2124
rect 7804 2096 7812 2104
rect 7772 2076 7780 2084
rect 7804 2076 7812 2084
rect 7804 1996 7812 2004
rect 7724 1936 7732 1944
rect 7500 1916 7508 1924
rect 7484 1896 7492 1904
rect 7532 1896 7540 1904
rect 7740 1896 7748 1904
rect 7772 1896 7780 1904
rect 7916 2556 7924 2564
rect 7884 2536 7892 2544
rect 8060 3096 8068 3104
rect 8060 3076 8068 3084
rect 8108 3296 8116 3304
rect 8092 3276 8100 3284
rect 8140 4156 8148 4164
rect 8140 4116 8148 4124
rect 8156 3716 8164 3724
rect 8156 3336 8164 3344
rect 8140 3096 8148 3104
rect 8060 2716 8068 2724
rect 8092 2676 8100 2684
rect 8108 2596 8116 2604
rect 8076 2576 8084 2584
rect 8108 2576 8116 2584
rect 7884 2336 7892 2344
rect 7916 2296 7924 2304
rect 7980 2302 7988 2304
rect 7980 2296 7988 2302
rect 7916 2276 7924 2284
rect 8108 2276 8116 2284
rect 7948 2136 7956 2144
rect 7836 2116 7844 2124
rect 7852 2116 7860 2124
rect 7868 2116 7876 2124
rect 7836 2096 7844 2104
rect 7836 1916 7844 1924
rect 7868 2096 7876 2104
rect 8060 2096 8068 2104
rect 7932 2076 7940 2084
rect 7964 1976 7972 1984
rect 8076 1936 8084 1944
rect 7868 1916 7876 1924
rect 7948 1916 7956 1924
rect 8060 1916 8068 1924
rect 7852 1896 7860 1904
rect 8012 1896 8020 1904
rect 7516 1876 7524 1884
rect 7596 1876 7604 1884
rect 7820 1876 7828 1884
rect 7852 1876 7860 1884
rect 7404 1776 7412 1784
rect 7564 1776 7572 1784
rect 7372 1756 7380 1764
rect 7340 1716 7348 1724
rect 7436 1718 7444 1724
rect 7436 1716 7444 1718
rect 7308 1696 7316 1704
rect 7356 1696 7364 1704
rect 7228 1676 7236 1684
rect 7436 1676 7444 1684
rect 7212 1656 7220 1664
rect 7148 1636 7156 1644
rect 7180 1636 7188 1644
rect 7404 1636 7412 1644
rect 6732 1576 6740 1584
rect 7004 1576 7012 1584
rect 7052 1576 7060 1584
rect 7100 1576 7108 1584
rect 6940 1556 6948 1564
rect 6860 1536 6868 1544
rect 6988 1536 6996 1544
rect 6748 1516 6756 1524
rect 6780 1516 6788 1524
rect 6860 1496 6868 1504
rect 6780 1476 6788 1484
rect 6828 1476 6836 1484
rect 6876 1476 6884 1484
rect 6812 1456 6820 1464
rect 6684 1436 6692 1444
rect 6748 1416 6756 1424
rect 6668 1396 6676 1404
rect 6588 1356 6596 1364
rect 6684 1336 6692 1344
rect 6556 1316 6564 1324
rect 6476 1276 6484 1284
rect 6348 1236 6356 1244
rect 6428 1236 6436 1244
rect 6316 1136 6324 1144
rect 6636 1276 6644 1284
rect 6588 1256 6596 1264
rect 6620 1256 6628 1264
rect 6556 1176 6564 1184
rect 6476 1116 6484 1124
rect 6508 1116 6516 1124
rect 6444 1096 6452 1104
rect 6572 1096 6580 1104
rect 6364 1076 6372 1084
rect 6332 1056 6340 1064
rect 6316 1036 6324 1044
rect 6348 1036 6356 1044
rect 6300 1016 6308 1024
rect 6300 956 6308 964
rect 6350 1006 6358 1014
rect 6364 1006 6372 1014
rect 6378 1006 6386 1014
rect 6476 1036 6484 1044
rect 6444 956 6452 964
rect 6380 936 6388 944
rect 5804 918 5812 924
rect 5804 916 5812 918
rect 5868 916 5876 924
rect 5996 916 6004 924
rect 6156 916 6164 924
rect 6172 916 6180 924
rect 6236 916 6244 924
rect 6284 916 6292 924
rect 5868 896 5876 904
rect 5740 876 5748 884
rect 5932 876 5940 884
rect 6140 876 6148 884
rect 5932 816 5940 824
rect 5788 676 5796 684
rect 5740 656 5748 664
rect 5772 656 5780 664
rect 5836 656 5844 664
rect 5804 636 5812 644
rect 5804 616 5812 624
rect 6140 736 6148 744
rect 5948 716 5956 724
rect 5980 716 5988 724
rect 5900 656 5908 664
rect 5772 576 5780 584
rect 5868 616 5876 624
rect 6012 696 6020 704
rect 6172 896 6180 904
rect 6284 896 6292 904
rect 6620 1236 6628 1244
rect 6668 1236 6676 1244
rect 6604 1136 6612 1144
rect 6652 1116 6660 1124
rect 6620 1076 6628 1084
rect 6588 1016 6596 1024
rect 6476 936 6484 944
rect 6796 1316 6804 1324
rect 6700 1236 6708 1244
rect 6780 1196 6788 1204
rect 6748 1176 6756 1184
rect 6764 1136 6772 1144
rect 6972 1476 6980 1484
rect 6908 1456 6916 1464
rect 6908 1336 6916 1344
rect 6828 1276 6836 1284
rect 6892 1276 6900 1284
rect 6812 1236 6820 1244
rect 6732 1096 6740 1104
rect 6652 936 6660 944
rect 6444 896 6452 904
rect 6700 936 6708 944
rect 6652 916 6660 924
rect 6796 1116 6804 1124
rect 6956 1276 6964 1284
rect 6924 1256 6932 1264
rect 7084 1556 7092 1564
rect 7196 1596 7204 1604
rect 7084 1496 7092 1504
rect 7196 1496 7204 1504
rect 7260 1496 7268 1504
rect 7052 1396 7060 1404
rect 7116 1396 7124 1404
rect 7292 1476 7300 1484
rect 7196 1416 7204 1424
rect 7100 1316 7108 1324
rect 7180 1316 7188 1324
rect 6988 1296 6996 1304
rect 7100 1296 7108 1304
rect 7084 1236 7092 1244
rect 6972 1216 6980 1224
rect 6860 1136 6868 1144
rect 6924 1136 6932 1144
rect 6812 1036 6820 1044
rect 7308 1396 7316 1404
rect 8012 1876 8020 1884
rect 7996 1856 8004 1864
rect 8044 1856 8052 1864
rect 7916 1776 7924 1784
rect 7948 1776 7956 1784
rect 7980 1756 7988 1764
rect 8012 1756 8020 1764
rect 7884 1736 7892 1744
rect 7980 1736 7988 1744
rect 7580 1656 7588 1664
rect 7500 1516 7508 1524
rect 7548 1516 7556 1524
rect 7484 1496 7492 1504
rect 7468 1476 7476 1484
rect 7644 1636 7652 1644
rect 7724 1536 7732 1544
rect 7772 1536 7780 1544
rect 7804 1536 7812 1544
rect 7900 1536 7908 1544
rect 7628 1516 7636 1524
rect 7692 1516 7700 1524
rect 7820 1516 7828 1524
rect 7868 1516 7876 1524
rect 7932 1516 7940 1524
rect 7964 1516 7972 1524
rect 7580 1496 7588 1504
rect 7596 1476 7604 1484
rect 7660 1476 7668 1484
rect 7580 1456 7588 1464
rect 7532 1376 7540 1384
rect 7404 1336 7412 1344
rect 7532 1336 7540 1344
rect 7676 1436 7684 1444
rect 7740 1476 7748 1484
rect 7724 1456 7732 1464
rect 7708 1416 7716 1424
rect 7356 1316 7364 1324
rect 7532 1316 7540 1324
rect 7628 1316 7636 1324
rect 7692 1316 7700 1324
rect 7628 1296 7636 1304
rect 7708 1296 7716 1304
rect 7244 1276 7252 1284
rect 7340 1276 7348 1284
rect 7516 1276 7524 1284
rect 7644 1276 7652 1284
rect 7244 1196 7252 1204
rect 7212 1136 7220 1144
rect 6956 1116 6964 1124
rect 7180 1116 7188 1124
rect 7244 1116 7252 1124
rect 6924 1076 6932 1084
rect 7132 1076 7140 1084
rect 6876 1036 6884 1044
rect 6844 1016 6852 1024
rect 6908 1016 6916 1024
rect 7036 1016 7044 1024
rect 7148 1036 7156 1044
rect 7132 976 7140 984
rect 7276 1076 7284 1084
rect 7708 1156 7716 1164
rect 7516 1136 7524 1144
rect 7596 1136 7604 1144
rect 7612 1136 7620 1144
rect 7644 1136 7652 1144
rect 7436 1116 7444 1124
rect 7372 1096 7380 1104
rect 7548 1096 7556 1104
rect 7324 1076 7332 1084
rect 7356 1076 7364 1084
rect 7372 1076 7380 1084
rect 7452 1076 7460 1084
rect 7484 1076 7492 1084
rect 7532 1076 7540 1084
rect 7420 1056 7428 1064
rect 7356 1036 7364 1044
rect 7308 1016 7316 1024
rect 7276 996 7284 1004
rect 6892 956 6900 964
rect 6924 956 6932 964
rect 7196 956 7204 964
rect 6972 936 6980 944
rect 6764 918 6772 924
rect 6764 916 6772 918
rect 6652 896 6660 904
rect 6732 896 6740 904
rect 6540 876 6548 884
rect 6604 876 6612 884
rect 6940 856 6948 864
rect 7372 936 7380 944
rect 7404 936 7412 944
rect 7068 916 7076 924
rect 7052 896 7060 904
rect 7404 916 7412 924
rect 7308 896 7316 904
rect 7244 856 7252 864
rect 7116 756 7124 764
rect 7212 756 7220 764
rect 6428 736 6436 744
rect 6492 736 6500 744
rect 6748 736 6756 744
rect 7004 736 7012 744
rect 7180 736 7188 744
rect 6396 716 6404 724
rect 6188 696 6196 704
rect 6332 696 6340 704
rect 6444 696 6452 704
rect 5948 576 5956 584
rect 5836 556 5844 564
rect 5932 556 5940 564
rect 5740 536 5748 544
rect 5820 536 5828 544
rect 5852 536 5860 544
rect 5676 516 5684 524
rect 5660 496 5668 504
rect 5548 296 5556 304
rect 5660 336 5668 344
rect 5596 316 5604 324
rect 5788 516 5796 524
rect 5692 456 5700 464
rect 5724 456 5732 464
rect 5740 336 5748 344
rect 5676 316 5684 324
rect 5772 316 5780 324
rect 5916 456 5924 464
rect 5804 316 5812 324
rect 5836 316 5844 324
rect 5900 316 5908 324
rect 5628 296 5636 304
rect 5692 296 5700 304
rect 5724 296 5732 304
rect 5628 256 5636 264
rect 5612 236 5620 244
rect 5564 156 5572 164
rect 6060 636 6068 644
rect 6012 536 6020 544
rect 6524 696 6532 704
rect 6476 676 6484 684
rect 6412 656 6420 664
rect 6268 636 6276 644
rect 6316 636 6324 644
rect 6350 606 6358 614
rect 6364 606 6372 614
rect 6378 606 6386 614
rect 6092 556 6100 564
rect 6236 556 6244 564
rect 6076 516 6084 524
rect 5948 296 5956 304
rect 5852 256 5860 264
rect 5708 236 5716 244
rect 5788 236 5796 244
rect 5772 176 5780 184
rect 6044 476 6052 484
rect 6124 476 6132 484
rect 6156 476 6164 484
rect 6284 576 6292 584
rect 6220 536 6228 544
rect 6316 556 6324 564
rect 6332 556 6340 564
rect 6444 556 6452 564
rect 6220 496 6228 504
rect 6188 416 6196 424
rect 5980 356 5988 364
rect 6412 536 6420 544
rect 6396 516 6404 524
rect 6412 496 6420 504
rect 6508 576 6516 584
rect 6508 556 6516 564
rect 6620 696 6628 704
rect 6652 696 6660 704
rect 6732 676 6740 684
rect 6556 576 6564 584
rect 6540 556 6548 564
rect 6524 536 6532 544
rect 6572 536 6580 544
rect 6940 716 6948 724
rect 6780 696 6788 704
rect 6812 696 6820 704
rect 6876 702 6884 704
rect 6876 696 6884 702
rect 6812 616 6820 624
rect 6684 576 6692 584
rect 6716 576 6724 584
rect 6764 576 6772 584
rect 6604 536 6612 544
rect 6812 536 6820 544
rect 6588 516 6596 524
rect 6748 516 6756 524
rect 6668 496 6676 504
rect 6476 476 6484 484
rect 6668 476 6676 484
rect 6716 476 6724 484
rect 6796 496 6804 504
rect 6508 456 6516 464
rect 6732 456 6740 464
rect 6300 396 6308 404
rect 6396 396 6404 404
rect 6284 376 6292 384
rect 6444 376 6452 384
rect 6812 376 6820 384
rect 6716 356 6724 364
rect 6236 296 6244 304
rect 6460 296 6468 304
rect 6524 302 6532 304
rect 6524 296 6532 302
rect 6700 296 6708 304
rect 6860 616 6868 624
rect 7116 696 7124 704
rect 7164 696 7172 704
rect 7244 696 7252 704
rect 7052 676 7060 684
rect 7276 676 7284 684
rect 7068 656 7076 664
rect 7132 656 7140 664
rect 7260 656 7268 664
rect 7020 576 7028 584
rect 6940 556 6948 564
rect 7276 596 7284 604
rect 7340 876 7348 884
rect 7388 876 7396 884
rect 7372 836 7380 844
rect 7372 716 7380 724
rect 7436 1036 7444 1044
rect 7436 976 7444 984
rect 7500 1056 7508 1064
rect 7548 1016 7556 1024
rect 7516 936 7524 944
rect 7484 916 7492 924
rect 7564 976 7572 984
rect 7660 1116 7668 1124
rect 7676 1096 7684 1104
rect 7580 916 7588 924
rect 7468 876 7476 884
rect 7500 876 7508 884
rect 7484 856 7492 864
rect 7420 756 7428 764
rect 7484 716 7492 724
rect 7516 716 7524 724
rect 7420 696 7428 704
rect 7324 676 7332 684
rect 7372 676 7380 684
rect 7404 676 7412 684
rect 7452 676 7460 684
rect 7548 676 7556 684
rect 7468 656 7476 664
rect 7644 936 7652 944
rect 7628 876 7636 884
rect 7612 836 7620 844
rect 7596 716 7604 724
rect 7756 1456 7764 1464
rect 7804 1456 7812 1464
rect 7772 1436 7780 1444
rect 7756 1416 7764 1424
rect 7852 1476 7860 1484
rect 7884 1476 7892 1484
rect 7820 1356 7828 1364
rect 7964 1456 7972 1464
rect 7900 1436 7908 1444
rect 7932 1436 7940 1444
rect 7948 1436 7956 1444
rect 7900 1356 7908 1364
rect 7836 1316 7844 1324
rect 7916 1316 7924 1324
rect 7996 1496 8004 1504
rect 8108 1496 8116 1504
rect 8012 1476 8020 1484
rect 8044 1456 8052 1464
rect 8028 1376 8036 1384
rect 7948 1336 7956 1344
rect 7756 1296 7764 1304
rect 7932 1296 7940 1304
rect 7772 1276 7780 1284
rect 7756 1096 7764 1104
rect 7884 1276 7892 1284
rect 7948 1276 7956 1284
rect 8012 1318 8020 1324
rect 8012 1316 8020 1318
rect 7980 1196 7988 1204
rect 8012 1196 8020 1204
rect 7980 1136 7988 1144
rect 7868 1096 7876 1104
rect 7900 1096 7908 1104
rect 7836 1076 7844 1084
rect 7868 1076 7876 1084
rect 7692 1056 7700 1064
rect 7724 1056 7732 1064
rect 7820 1056 7828 1064
rect 7852 1056 7860 1064
rect 7964 1056 7972 1064
rect 7708 976 7716 984
rect 7788 1016 7796 1024
rect 7740 996 7748 1004
rect 7740 956 7748 964
rect 7804 936 7812 944
rect 7724 916 7732 924
rect 7900 976 7908 984
rect 7852 916 7860 924
rect 7884 916 7892 924
rect 8044 1336 8052 1344
rect 8060 1156 8068 1164
rect 8108 1056 8116 1064
rect 8060 1016 8068 1024
rect 8092 1016 8100 1024
rect 8012 956 8020 964
rect 8108 976 8116 984
rect 8156 2896 8164 2904
rect 8156 2096 8164 2104
rect 8156 1936 8164 1944
rect 8140 1916 8148 1924
rect 8140 1156 8148 1164
rect 7740 896 7748 904
rect 7852 896 7860 904
rect 7884 896 7892 904
rect 7996 896 8004 904
rect 7756 836 7764 844
rect 7804 716 7812 724
rect 7852 716 7860 724
rect 7788 696 7796 704
rect 7772 676 7780 684
rect 7724 656 7732 664
rect 7276 576 7284 584
rect 7308 576 7316 584
rect 7260 556 7268 564
rect 7020 536 7028 544
rect 7084 536 7092 544
rect 6860 516 6868 524
rect 7036 516 7044 524
rect 7084 516 7092 524
rect 7004 496 7012 504
rect 6988 476 6996 484
rect 6956 356 6964 364
rect 7020 356 7028 364
rect 6892 336 6900 344
rect 6924 336 6932 344
rect 6012 276 6020 284
rect 6108 276 6116 284
rect 6556 276 6564 284
rect 6652 276 6660 284
rect 6844 276 6852 284
rect 6892 276 6900 284
rect 5980 236 5988 244
rect 5756 156 5764 164
rect 5852 156 5860 164
rect 5932 156 5940 164
rect 5964 156 5972 164
rect 5260 136 5268 144
rect 5324 136 5332 144
rect 5468 136 5476 144
rect 5580 136 5588 144
rect 5708 136 5716 144
rect 5964 116 5972 124
rect 6092 196 6100 204
rect 6252 196 6260 204
rect 6108 156 6116 164
rect 6236 156 6244 164
rect 6284 156 6292 164
rect 3692 96 3700 104
rect 3772 96 3780 104
rect 3868 96 3876 104
rect 4092 96 4100 104
rect 4284 96 4292 104
rect 4396 96 4404 104
rect 4460 96 4468 104
rect 4700 96 4708 104
rect 4748 96 4756 104
rect 4828 96 4836 104
rect 4924 96 4932 104
rect 5052 96 5060 104
rect 5148 96 5156 104
rect 5244 96 5252 104
rect 5356 96 5364 104
rect 5660 96 5668 104
rect 5724 96 5732 104
rect 5756 96 5764 104
rect 5884 96 5892 104
rect 6012 96 6020 104
rect 6620 256 6628 264
rect 6796 256 6804 264
rect 6588 236 6596 244
rect 6350 206 6358 214
rect 6364 206 6372 214
rect 6378 206 6386 214
rect 6588 156 6596 164
rect 6604 156 6612 164
rect 6476 140 6484 144
rect 6476 136 6484 140
rect 6524 136 6532 144
rect 6540 136 6548 144
rect 6572 136 6580 144
rect 6396 116 6404 124
rect 6716 196 6724 204
rect 6780 196 6788 204
rect 6652 176 6660 184
rect 6636 136 6644 144
rect 6668 156 6676 164
rect 6876 256 6884 264
rect 6844 236 6852 244
rect 6860 236 6868 244
rect 6732 176 6740 184
rect 6812 176 6820 184
rect 6812 156 6820 164
rect 6780 136 6788 144
rect 6844 136 6852 144
rect 7052 476 7060 484
rect 6972 276 6980 284
rect 6988 256 6996 264
rect 7004 236 7012 244
rect 6924 216 6932 224
rect 6956 216 6964 224
rect 6668 116 6676 124
rect 6764 116 6772 124
rect 6796 116 6804 124
rect 6892 116 6900 124
rect 6988 196 6996 204
rect 7084 356 7092 364
rect 7372 596 7380 604
rect 7180 496 7188 504
rect 7132 356 7140 364
rect 7116 336 7124 344
rect 7196 336 7204 344
rect 7148 316 7156 324
rect 7132 296 7140 304
rect 7244 316 7252 324
rect 7228 296 7236 304
rect 7052 276 7060 284
rect 7036 256 7044 264
rect 7100 256 7108 264
rect 7260 296 7268 304
rect 7324 302 7332 304
rect 7324 296 7332 302
rect 7212 216 7220 224
rect 7020 196 7028 204
rect 7484 576 7492 584
rect 7516 576 7524 584
rect 7436 536 7444 544
rect 7452 376 7460 384
rect 7676 556 7684 564
rect 7580 536 7588 544
rect 7532 516 7540 524
rect 7628 516 7636 524
rect 7772 516 7780 524
rect 7788 396 7796 404
rect 7500 316 7508 324
rect 7708 316 7716 324
rect 7692 296 7700 304
rect 7740 296 7748 304
rect 7468 276 7476 284
rect 7660 276 7668 284
rect 7708 276 7716 284
rect 7740 276 7748 284
rect 7628 236 7636 244
rect 7276 156 7284 164
rect 7340 156 7348 164
rect 7532 156 7540 164
rect 7116 136 7124 144
rect 7308 136 7316 144
rect 7404 136 7412 144
rect 8076 736 8084 744
rect 7980 716 7988 724
rect 8060 716 8068 724
rect 7900 696 7908 704
rect 8012 696 8020 704
rect 7836 676 7844 684
rect 7868 676 7876 684
rect 7980 676 7988 684
rect 7804 296 7812 304
rect 7836 636 7844 644
rect 7852 396 7860 404
rect 7996 656 8004 664
rect 7964 636 7972 644
rect 7916 616 7924 624
rect 7964 516 7972 524
rect 7980 516 7988 524
rect 8028 656 8036 664
rect 8012 616 8020 624
rect 8060 616 8068 624
rect 8108 716 8116 724
rect 8092 696 8100 704
rect 8108 676 8116 684
rect 8092 656 8100 664
rect 8156 656 8164 664
rect 8140 636 8148 644
rect 8028 516 8036 524
rect 8044 516 8052 524
rect 8060 496 8068 504
rect 8124 496 8132 504
rect 8092 476 8100 484
rect 7916 396 7924 404
rect 7884 316 7892 324
rect 7916 316 7924 324
rect 7820 276 7828 284
rect 7852 216 7860 224
rect 7868 196 7876 204
rect 7756 176 7764 184
rect 7836 176 7844 184
rect 7852 156 7860 164
rect 8108 396 8116 404
rect 7932 296 7940 304
rect 7980 296 7988 304
rect 8060 296 8068 304
rect 7996 276 8004 284
rect 7916 196 7924 204
rect 7868 136 7876 144
rect 6940 116 6948 124
rect 6972 116 6980 124
rect 7052 116 7060 124
rect 7356 116 7364 124
rect 7420 116 7428 124
rect 7596 118 7604 124
rect 7596 116 7604 118
rect 7932 136 7940 144
rect 8028 276 8036 284
rect 8012 236 8020 244
rect 7964 216 7972 224
rect 7996 176 8004 184
rect 7964 156 7972 164
rect 8012 156 8020 164
rect 7932 116 7940 124
rect 8092 256 8100 264
rect 8092 236 8100 244
rect 8076 156 8084 164
rect 8060 136 8068 144
rect 8092 136 8100 144
rect 8060 116 8068 124
rect 6460 96 6468 104
rect 6620 96 6628 104
rect 6748 96 6756 104
rect 6924 96 6932 104
rect 7020 96 7028 104
rect 7052 96 7060 104
rect 7228 96 7236 104
rect 7388 96 7396 104
rect 7420 96 7428 104
rect 8028 96 8036 104
rect 8076 96 8084 104
rect 8156 296 8164 304
rect 2060 76 2068 84
rect 6204 76 6212 84
rect 6316 76 6324 84
rect 7356 76 7364 84
rect 1742 6 1750 14
rect 1756 6 1764 14
rect 1770 6 1778 14
rect 4814 6 4822 14
rect 4828 6 4836 14
rect 4842 6 4850 14
<< metal3 >>
rect 3272 5814 3320 5816
rect 3272 5806 3276 5814
rect 3286 5806 3292 5814
rect 3300 5806 3306 5814
rect 3316 5806 3320 5814
rect 3272 5804 3320 5806
rect 6344 5814 6392 5816
rect 6344 5806 6348 5814
rect 6358 5806 6364 5814
rect 6372 5806 6378 5814
rect 6388 5806 6392 5814
rect 6344 5804 6392 5806
rect 2820 5797 2844 5803
rect 3028 5797 3068 5803
rect 3620 5797 3644 5803
rect 6164 5797 6204 5803
rect 2740 5777 2828 5783
rect 3156 5777 3292 5783
rect 4516 5777 4764 5783
rect 4772 5777 5020 5783
rect 6148 5777 6204 5783
rect 692 5757 940 5763
rect 996 5757 1036 5763
rect 1044 5757 1116 5763
rect 1124 5757 1276 5763
rect 1284 5757 1484 5763
rect 2372 5757 2460 5763
rect 2468 5757 2588 5763
rect 3684 5757 3884 5763
rect 3956 5757 4156 5763
rect 4564 5757 4588 5763
rect 5044 5757 5452 5763
rect 5556 5757 5612 5763
rect 5844 5757 5884 5763
rect 6116 5757 6188 5763
rect 6196 5757 6572 5763
rect 6580 5757 6780 5763
rect 7060 5757 7324 5763
rect 292 5737 332 5743
rect 340 5737 636 5743
rect 884 5737 1148 5743
rect 1492 5737 1660 5743
rect 1668 5737 1868 5743
rect 1876 5737 2012 5743
rect 2020 5737 2204 5743
rect 2612 5737 2652 5743
rect 2996 5737 3356 5743
rect 3556 5737 3740 5743
rect 3876 5737 3964 5743
rect 4404 5737 4988 5743
rect 4996 5737 5084 5743
rect 5188 5737 5244 5743
rect 5492 5737 5612 5743
rect 5700 5737 5836 5743
rect 5908 5737 6092 5743
rect 6372 5737 6444 5743
rect 6452 5737 6652 5743
rect 6660 5737 6908 5743
rect 7124 5737 7164 5743
rect 7348 5737 7356 5743
rect 7620 5737 7644 5743
rect 7876 5737 7964 5743
rect 7972 5737 7996 5743
rect 100 5717 204 5723
rect 244 5717 380 5723
rect 516 5717 700 5723
rect 932 5717 1004 5723
rect 1012 5717 1036 5723
rect 1044 5717 1116 5723
rect 1124 5717 1164 5723
rect 1332 5717 1420 5723
rect 1796 5717 1820 5723
rect 2068 5717 2252 5723
rect 2276 5717 2380 5723
rect 2580 5717 2700 5723
rect 2820 5717 2924 5723
rect 3284 5717 3404 5723
rect 3460 5717 3596 5723
rect 3604 5717 3676 5723
rect 4100 5717 4284 5723
rect 4468 5717 4524 5723
rect 4564 5717 4620 5723
rect 4692 5717 4844 5723
rect 5076 5717 5132 5723
rect 5188 5717 5500 5723
rect 5620 5717 5692 5723
rect 5700 5717 5772 5723
rect 5780 5717 5820 5723
rect 5844 5717 5980 5723
rect 6084 5717 6316 5723
rect 6724 5717 6748 5723
rect 7108 5717 7132 5723
rect 7156 5717 7324 5723
rect 132 5697 556 5703
rect 564 5697 748 5703
rect 1204 5697 1276 5703
rect 1284 5697 1420 5703
rect 1588 5697 1644 5703
rect 1684 5697 1724 5703
rect 1796 5697 2332 5703
rect 2388 5697 2492 5703
rect 2628 5697 2812 5703
rect 3044 5697 3228 5703
rect 3540 5697 3724 5703
rect 3732 5697 3772 5703
rect 3780 5697 4060 5703
rect 4068 5697 4108 5703
rect 4845 5703 4851 5716
rect 4845 5697 5212 5703
rect 5380 5697 5516 5703
rect 5668 5697 5788 5703
rect 5812 5697 5852 5703
rect 6948 5697 7004 5703
rect 7028 5697 7084 5703
rect 7204 5697 7260 5703
rect 372 5677 428 5683
rect 436 5677 540 5683
rect 916 5677 1100 5683
rect 1108 5677 1180 5683
rect 1252 5677 1324 5683
rect 1364 5677 1468 5683
rect 1700 5677 1900 5683
rect 2420 5677 2476 5683
rect 2484 5677 2636 5683
rect 2644 5677 2716 5683
rect 2724 5677 2780 5683
rect 2788 5677 3052 5683
rect 3060 5677 3196 5683
rect 3204 5677 3532 5683
rect 3636 5677 3836 5683
rect 3844 5677 3996 5683
rect 4004 5677 4492 5683
rect 4516 5677 4988 5683
rect 5124 5677 5388 5683
rect 5492 5677 5692 5683
rect 5716 5677 5772 5683
rect 5789 5683 5795 5696
rect 5789 5677 5868 5683
rect 5876 5677 5884 5683
rect 5924 5677 6092 5683
rect 6964 5677 7132 5683
rect 7156 5677 7212 5683
rect 212 5657 364 5663
rect 724 5657 1020 5663
rect 1124 5657 1340 5663
rect 1620 5657 1788 5663
rect 1828 5657 1980 5663
rect 1988 5657 2444 5663
rect 2548 5657 2668 5663
rect 2676 5657 2828 5663
rect 2836 5657 3084 5663
rect 3092 5657 3628 5663
rect 5012 5657 5052 5663
rect 5060 5657 5468 5663
rect 5572 5657 5756 5663
rect 5844 5657 6060 5663
rect 6980 5657 7100 5663
rect 7108 5657 7212 5663
rect 1556 5637 1564 5643
rect 1844 5637 1884 5643
rect 4004 5637 4044 5643
rect 4340 5637 4620 5643
rect 5428 5637 5532 5643
rect 5812 5637 5884 5643
rect 5892 5637 5948 5643
rect 6996 5637 7276 5643
rect 7716 5637 8012 5643
rect 4020 5617 4204 5623
rect 5732 5617 5996 5623
rect 7460 5617 7836 5623
rect 1736 5614 1784 5616
rect 1736 5606 1740 5614
rect 1750 5606 1756 5614
rect 1764 5606 1770 5614
rect 1780 5606 1784 5614
rect 1736 5604 1784 5606
rect 4808 5614 4856 5616
rect 4808 5606 4812 5614
rect 4822 5606 4828 5614
rect 4836 5606 4842 5614
rect 4852 5606 4856 5614
rect 4808 5604 4856 5606
rect 916 5597 956 5603
rect 3092 5597 3148 5603
rect 3908 5597 4092 5603
rect 4116 5597 4172 5603
rect 4276 5597 4380 5603
rect 5636 5597 5740 5603
rect 5764 5597 5916 5603
rect 84 5577 492 5583
rect 1604 5577 1980 5583
rect 2708 5577 2796 5583
rect 2804 5577 3116 5583
rect 3124 5577 3596 5583
rect 3604 5577 3964 5583
rect 3972 5577 4108 5583
rect 4740 5577 4972 5583
rect 5396 5577 5580 5583
rect 5588 5577 5740 5583
rect 5748 5577 6188 5583
rect 7412 5577 7420 5583
rect 404 5557 444 5563
rect 996 5557 1244 5563
rect 1636 5557 1932 5563
rect 4388 5557 4412 5563
rect 4596 5557 4812 5563
rect 4980 5557 5564 5563
rect 5812 5557 5900 5563
rect 7892 5557 7948 5563
rect 1076 5537 1100 5543
rect 1188 5537 1372 5543
rect 1572 5537 1612 5543
rect 1860 5537 1996 5543
rect 2004 5537 2028 5543
rect 2036 5537 2092 5543
rect 2164 5537 2220 5543
rect 2676 5537 2908 5543
rect 4404 5537 4572 5543
rect 5028 5537 5052 5543
rect 5108 5537 5164 5543
rect 5780 5537 5836 5543
rect 6212 5537 6508 5543
rect 6516 5537 6700 5543
rect 6900 5537 7420 5543
rect 7764 5537 7868 5543
rect 7924 5537 7996 5543
rect 260 5517 300 5523
rect 516 5517 556 5523
rect 980 5517 1148 5523
rect 1156 5517 1228 5523
rect 1236 5517 1340 5523
rect 2036 5517 2204 5523
rect 2212 5517 2348 5523
rect 2548 5517 2860 5523
rect 3444 5517 3548 5523
rect 4132 5517 4332 5523
rect 4340 5517 4380 5523
rect 4532 5517 4556 5523
rect 4980 5517 5068 5523
rect 5876 5517 6028 5523
rect 6036 5517 6140 5523
rect 6596 5517 6620 5523
rect 6628 5517 6684 5523
rect 7172 5517 7468 5523
rect 7604 5517 7852 5523
rect 7860 5517 8076 5523
rect 212 5497 332 5503
rect 372 5497 428 5503
rect 436 5497 572 5503
rect 980 5497 1052 5503
rect 1364 5497 1436 5503
rect 1940 5497 1980 5503
rect 2228 5497 2252 5503
rect 2484 5497 2492 5503
rect 2676 5497 2844 5503
rect 2948 5497 3004 5503
rect 3332 5497 3436 5503
rect 3476 5497 3532 5503
rect 3572 5497 3644 5503
rect 3780 5497 3916 5503
rect 3988 5497 4044 5503
rect 4228 5497 4364 5503
rect 4372 5497 4444 5503
rect 4788 5497 4828 5503
rect 4836 5497 4940 5503
rect 5076 5497 5148 5503
rect 5188 5497 5388 5503
rect 5796 5497 5852 5503
rect 5892 5497 5900 5503
rect 6004 5497 6028 5503
rect 6548 5497 6572 5503
rect 6612 5497 6636 5503
rect 6692 5497 6780 5503
rect 7140 5497 7276 5503
rect 7876 5497 7900 5503
rect 8084 5497 8124 5503
rect 228 5477 300 5483
rect 356 5477 380 5483
rect 388 5477 412 5483
rect 484 5477 604 5483
rect 612 5477 764 5483
rect 1124 5477 1132 5483
rect 1236 5477 1452 5483
rect 1956 5477 2092 5483
rect 2100 5477 2124 5483
rect 2132 5477 2172 5483
rect 2452 5477 2492 5483
rect 2900 5477 3036 5483
rect 3428 5477 3516 5483
rect 3524 5477 3580 5483
rect 3924 5477 4076 5483
rect 4100 5477 4284 5483
rect 4292 5477 4540 5483
rect 4548 5477 4620 5483
rect 4804 5477 5132 5483
rect 5524 5477 5676 5483
rect 5684 5477 5756 5483
rect 5764 5477 6044 5483
rect 6052 5477 6252 5483
rect 6260 5477 6380 5483
rect 6388 5477 6492 5483
rect 6500 5477 6652 5483
rect 7124 5477 7228 5483
rect 7236 5477 7260 5483
rect 7524 5477 7692 5483
rect 7828 5477 7996 5483
rect 8116 5477 8124 5483
rect 196 5457 316 5463
rect 404 5457 428 5463
rect 900 5457 940 5463
rect 948 5457 1052 5463
rect 1060 5457 1132 5463
rect 1172 5457 1292 5463
rect 1556 5457 1644 5463
rect 1764 5457 1868 5463
rect 1876 5457 1996 5463
rect 2148 5457 2300 5463
rect 2948 5457 3100 5463
rect 3636 5457 3708 5463
rect 4260 5457 4316 5463
rect 4324 5457 4332 5463
rect 4340 5457 4460 5463
rect 4468 5457 4556 5463
rect 4900 5457 5084 5463
rect 5092 5457 5116 5463
rect 5124 5457 5212 5463
rect 5236 5457 5276 5463
rect 5444 5457 5580 5463
rect 5892 5457 6108 5463
rect 6116 5457 6716 5463
rect 6884 5457 7084 5463
rect 7092 5457 7116 5463
rect 7188 5457 7548 5463
rect 7844 5457 7948 5463
rect 276 5437 396 5443
rect 468 5437 620 5443
rect 628 5437 876 5443
rect 1044 5437 1404 5443
rect 1908 5437 1964 5443
rect 1972 5437 2300 5443
rect 2308 5437 5244 5443
rect 5556 5437 5708 5443
rect 5716 5437 5932 5443
rect 5940 5437 5948 5443
rect 6388 5437 6428 5443
rect 6708 5437 6748 5443
rect 7044 5437 7068 5443
rect 7076 5437 7340 5443
rect 7348 5437 7420 5443
rect 7636 5437 7692 5443
rect 7700 5437 8044 5443
rect 852 5417 972 5423
rect 1028 5417 1212 5423
rect 1812 5417 2028 5423
rect 3140 5417 3228 5423
rect 3716 5417 3836 5423
rect 4180 5417 4332 5423
rect 4340 5417 4492 5423
rect 4740 5417 4748 5423
rect 4980 5417 5020 5423
rect 5028 5417 5068 5423
rect 5076 5417 5148 5423
rect 5156 5417 5196 5423
rect 5908 5417 6188 5423
rect 7956 5417 7996 5423
rect 3272 5414 3320 5416
rect 3272 5406 3276 5414
rect 3286 5406 3292 5414
rect 3300 5406 3306 5414
rect 3316 5406 3320 5414
rect 3272 5404 3320 5406
rect 6344 5414 6392 5416
rect 6344 5406 6348 5414
rect 6358 5406 6364 5414
rect 6372 5406 6378 5414
rect 6388 5406 6392 5414
rect 6344 5404 6392 5406
rect 420 5397 540 5403
rect 548 5397 851 5403
rect 845 5384 851 5397
rect 1220 5397 1260 5403
rect 1268 5397 1308 5403
rect 1668 5397 1820 5403
rect 2052 5397 2380 5403
rect 2772 5397 2828 5403
rect 4020 5397 4060 5403
rect 4068 5397 4268 5403
rect 6724 5397 6796 5403
rect 7108 5397 7244 5403
rect 20 5377 28 5383
rect 36 5377 204 5383
rect 308 5377 556 5383
rect 580 5377 828 5383
rect 852 5377 924 5383
rect 932 5377 1100 5383
rect 1108 5377 1148 5383
rect 1284 5377 1308 5383
rect 1652 5377 2044 5383
rect 2852 5377 3500 5383
rect 4212 5377 4300 5383
rect 4932 5377 5004 5383
rect 5012 5377 5100 5383
rect 5108 5377 5116 5383
rect 6052 5377 6284 5383
rect 6372 5377 6588 5383
rect 6772 5377 7132 5383
rect 7284 5377 7404 5383
rect 7460 5377 7772 5383
rect 8036 5377 8076 5383
rect 324 5357 364 5363
rect 372 5357 460 5363
rect 564 5357 636 5363
rect 660 5357 700 5363
rect 708 5357 940 5363
rect 948 5357 1692 5363
rect 1700 5357 1740 5363
rect 2036 5357 2204 5363
rect 2420 5357 2620 5363
rect 3108 5357 3132 5363
rect 3172 5357 3356 5363
rect 3524 5357 3772 5363
rect 3876 5357 3916 5363
rect 4036 5357 4316 5363
rect 5012 5357 5196 5363
rect 5220 5357 5340 5363
rect 5380 5357 6732 5363
rect 6740 5357 6780 5363
rect 7076 5357 7196 5363
rect 7972 5357 8140 5363
rect 228 5337 284 5343
rect 324 5337 396 5343
rect 628 5337 716 5343
rect 1684 5337 2092 5343
rect 2180 5337 2236 5343
rect 2292 5337 2444 5343
rect 2612 5337 2668 5343
rect 2676 5337 2908 5343
rect 2916 5337 3004 5343
rect 3012 5337 3052 5343
rect 3092 5337 3164 5343
rect 3540 5337 3580 5343
rect 3652 5337 3692 5343
rect 4100 5337 4156 5343
rect 4228 5337 4284 5343
rect 4292 5337 4348 5343
rect 4740 5337 4764 5343
rect 4996 5337 5020 5343
rect 5300 5337 5436 5343
rect 5508 5337 5548 5343
rect 5572 5337 6108 5343
rect 6148 5337 6220 5343
rect 6228 5337 6284 5343
rect 6292 5337 6316 5343
rect 6324 5337 6524 5343
rect 6532 5337 6588 5343
rect 6804 5337 7004 5343
rect 7028 5337 7084 5343
rect 7252 5337 7356 5343
rect 7716 5337 7836 5343
rect 7844 5337 7868 5343
rect 7876 5337 7932 5343
rect 7988 5337 8028 5343
rect 148 5317 252 5323
rect 276 5317 316 5323
rect 452 5317 540 5323
rect 548 5317 684 5323
rect 820 5317 844 5323
rect 916 5317 1244 5323
rect 1252 5317 1292 5323
rect 1380 5317 1500 5323
rect 1716 5317 1916 5323
rect 1988 5317 2028 5323
rect 2260 5317 2332 5323
rect 2388 5317 2476 5323
rect 2868 5317 2892 5323
rect 3076 5317 3180 5323
rect 3188 5317 3564 5323
rect 3572 5317 3676 5323
rect 3684 5317 3884 5323
rect 3892 5317 3948 5323
rect 3956 5317 4012 5323
rect 4148 5317 4172 5323
rect 4196 5317 4236 5323
rect 4436 5317 4492 5323
rect 4564 5317 4636 5323
rect 4740 5317 5132 5323
rect 5140 5317 5180 5323
rect 5188 5317 5228 5323
rect 5348 5317 5420 5323
rect 5444 5317 5484 5323
rect 5492 5317 5516 5323
rect 5668 5317 5692 5323
rect 5700 5317 5772 5323
rect 5780 5317 5996 5323
rect 6276 5317 6316 5323
rect 6340 5317 6460 5323
rect 6532 5317 6572 5323
rect 6580 5317 6700 5323
rect 6996 5317 7180 5323
rect 7300 5317 7388 5323
rect 7412 5317 7452 5323
rect 7764 5317 7900 5323
rect 7908 5317 7948 5323
rect 8004 5317 8044 5323
rect 8132 5317 8140 5323
rect 356 5297 460 5303
rect 468 5297 668 5303
rect 820 5297 860 5303
rect 1140 5297 1260 5303
rect 1300 5297 1356 5303
rect 2084 5297 2396 5303
rect 3060 5297 3324 5303
rect 3988 5297 4220 5303
rect 4276 5297 4380 5303
rect 4916 5297 5052 5303
rect 5204 5297 5244 5303
rect 5956 5297 6220 5303
rect 6388 5297 6476 5303
rect 6484 5297 6492 5303
rect 6548 5297 6620 5303
rect 6884 5297 7020 5303
rect 7108 5297 7324 5303
rect 7748 5297 7772 5303
rect 7796 5297 7820 5303
rect 7828 5297 7884 5303
rect 7892 5297 8028 5303
rect 436 5277 460 5283
rect 532 5277 556 5283
rect 676 5277 1756 5283
rect 2004 5277 2108 5283
rect 2116 5277 2268 5283
rect 2612 5277 2636 5283
rect 2644 5277 5340 5283
rect 6340 5277 6636 5283
rect 7156 5277 7228 5283
rect 7236 5277 7292 5283
rect 7812 5277 7852 5283
rect 7860 5277 7916 5283
rect 7924 5277 7980 5283
rect 7988 5277 8012 5283
rect 452 5257 652 5263
rect 2228 5257 2364 5263
rect 3220 5257 3484 5263
rect 3556 5257 3660 5263
rect 3668 5257 3980 5263
rect 4612 5257 4940 5263
rect 6036 5257 6172 5263
rect 6356 5257 6444 5263
rect 6452 5257 6540 5263
rect 7172 5257 7436 5263
rect 7572 5257 7772 5263
rect 1572 5237 4092 5243
rect 4452 5237 4780 5243
rect 6276 5237 6300 5243
rect 7684 5237 7820 5243
rect 7828 5237 7868 5243
rect 612 5217 1708 5223
rect 3028 5217 3116 5223
rect 3172 5217 3548 5223
rect 5844 5217 6828 5223
rect 1736 5214 1784 5216
rect 1736 5206 1740 5214
rect 1750 5206 1756 5214
rect 1764 5206 1770 5214
rect 1780 5206 1784 5214
rect 1736 5204 1784 5206
rect 4808 5214 4856 5216
rect 4808 5206 4812 5214
rect 4822 5206 4828 5214
rect 4836 5206 4842 5214
rect 4852 5206 4856 5214
rect 4808 5204 4856 5206
rect 1188 5197 1356 5203
rect 1364 5197 1612 5203
rect 3604 5197 3868 5203
rect 3876 5197 3900 5203
rect 6212 5197 6444 5203
rect 212 5177 2140 5183
rect 2356 5177 4828 5183
rect 4916 5177 5148 5183
rect 5284 5177 5836 5183
rect 5956 5177 6364 5183
rect 1316 5157 3804 5163
rect 4644 5157 4876 5163
rect 6212 5157 6236 5163
rect 6308 5157 6332 5163
rect 6468 5157 6508 5163
rect 6516 5157 6604 5163
rect 7140 5157 7164 5163
rect 7300 5157 7484 5163
rect 7812 5157 7852 5163
rect 1124 5137 1276 5143
rect 1284 5137 1308 5143
rect 2228 5137 2332 5143
rect 2548 5137 2748 5143
rect 2756 5137 2860 5143
rect 3220 5137 3516 5143
rect 3620 5137 3756 5143
rect 3796 5137 4012 5143
rect 4740 5137 4892 5143
rect 6244 5137 6348 5143
rect 6420 5137 6572 5143
rect 7172 5137 7388 5143
rect 7716 5137 7884 5143
rect 1924 5117 2188 5123
rect 2244 5117 2444 5123
rect 2452 5117 2460 5123
rect 2468 5117 2492 5123
rect 2564 5117 2620 5123
rect 2676 5117 2732 5123
rect 2932 5117 2956 5123
rect 3236 5117 3244 5123
rect 3364 5117 3516 5123
rect 3556 5117 3628 5123
rect 3732 5117 3788 5123
rect 3844 5117 3852 5123
rect 4148 5117 4204 5123
rect 4756 5117 4796 5123
rect 4932 5117 5020 5123
rect 5412 5117 5532 5123
rect 6148 5117 6524 5123
rect 7508 5117 7676 5123
rect 7860 5117 7900 5123
rect 7940 5117 8060 5123
rect 8084 5117 8092 5123
rect 84 5097 204 5103
rect 244 5097 268 5103
rect 500 5097 604 5103
rect 996 5097 1148 5103
rect 1316 5097 1372 5103
rect 2036 5097 2428 5103
rect 2436 5097 2572 5103
rect 2580 5097 2883 5103
rect 2877 5084 2883 5097
rect 3108 5097 3340 5103
rect 3476 5097 3612 5103
rect 3652 5097 3724 5103
rect 3908 5097 3980 5103
rect 4084 5097 4268 5103
rect 4276 5097 4476 5103
rect 4532 5097 4716 5103
rect 5044 5097 5164 5103
rect 5396 5097 5420 5103
rect 5428 5097 5452 5103
rect 5924 5097 6204 5103
rect 6228 5097 6428 5103
rect 6436 5097 6492 5103
rect 6900 5097 6908 5103
rect 7684 5097 7740 5103
rect 7844 5097 8044 5103
rect 8100 5097 8195 5103
rect 292 5077 364 5083
rect 1076 5077 1132 5083
rect 1412 5077 1468 5083
rect 1524 5077 1868 5083
rect 2164 5077 2236 5083
rect 2260 5077 2268 5083
rect 2276 5077 2476 5083
rect 2532 5077 2588 5083
rect 2612 5077 2668 5083
rect 2884 5077 3004 5083
rect 3220 5077 3372 5083
rect 3428 5077 3452 5083
rect 3556 5077 3580 5083
rect 3588 5077 3740 5083
rect 3892 5077 3932 5083
rect 4708 5077 4748 5083
rect 4804 5077 4972 5083
rect 5108 5077 5260 5083
rect 5444 5077 5500 5083
rect 5524 5077 5756 5083
rect 6180 5077 6300 5083
rect 6340 5077 6476 5083
rect 6548 5077 6732 5083
rect 6740 5077 6828 5083
rect 7076 5077 7228 5083
rect 7236 5077 7292 5083
rect 7508 5077 7692 5083
rect 7700 5077 7820 5083
rect 7860 5077 8028 5083
rect 132 5057 204 5063
rect 564 5057 588 5063
rect 1124 5057 1244 5063
rect 1252 5057 1308 5063
rect 1316 5057 1340 5063
rect 2148 5057 2188 5063
rect 2676 5057 2700 5063
rect 2964 5057 3004 5063
rect 3348 5057 3484 5063
rect 3508 5057 3580 5063
rect 3620 5057 3660 5063
rect 3844 5057 4140 5063
rect 4148 5057 4444 5063
rect 4452 5057 4652 5063
rect 4708 5057 4940 5063
rect 5236 5057 5308 5063
rect 5316 5057 5900 5063
rect 5908 5057 6956 5063
rect 6964 5057 7164 5063
rect 7172 5057 7196 5063
rect 7204 5057 7356 5063
rect 7412 5057 7740 5063
rect 7828 5057 8012 5063
rect 196 5037 524 5043
rect 1108 5037 1180 5043
rect 1236 5037 1356 5043
rect 3892 5037 3916 5043
rect 4196 5037 4412 5043
rect 4644 5037 4780 5043
rect 4884 5037 5500 5043
rect 5524 5037 5564 5043
rect 6164 5037 6380 5043
rect 6580 5037 6636 5043
rect 6740 5037 6764 5043
rect 6916 5037 7052 5043
rect 7220 5037 7244 5043
rect 7252 5037 7372 5043
rect 7492 5037 7820 5043
rect 3012 5017 3052 5023
rect 3876 5017 3900 5023
rect 5556 5017 5596 5023
rect 5796 5017 5996 5023
rect 6708 5017 6988 5023
rect 7332 5017 7404 5023
rect 7636 5017 7676 5023
rect 7732 5017 7980 5023
rect 3272 5014 3320 5016
rect 3272 5006 3276 5014
rect 3286 5006 3292 5014
rect 3300 5006 3306 5014
rect 3316 5006 3320 5014
rect 3272 5004 3320 5006
rect 6344 5014 6392 5016
rect 6344 5006 6348 5014
rect 6358 5006 6364 5014
rect 6372 5006 6378 5014
rect 6388 5006 6392 5014
rect 6344 5004 6392 5006
rect 212 4997 284 5003
rect 356 4997 460 5003
rect 1156 4997 1747 5003
rect 148 4977 396 4983
rect 644 4977 780 4983
rect 1268 4977 1548 4983
rect 1741 4983 1747 4997
rect 2308 4997 2572 5003
rect 2580 4997 2924 5003
rect 2932 4997 3212 5003
rect 3572 4997 3644 5003
rect 3652 4997 3692 5003
rect 4740 4997 4748 5003
rect 5524 4997 5772 5003
rect 7396 4997 7612 5003
rect 7780 4997 7948 5003
rect 1741 4977 2588 4983
rect 2596 4977 2876 4983
rect 2916 4977 3100 4983
rect 3108 4977 3228 4983
rect 3236 4977 3388 4983
rect 3748 4977 3820 4983
rect 3828 4977 3980 4983
rect 4788 4977 4908 4983
rect 5540 4977 5708 4983
rect 6292 4977 6764 4983
rect 7140 4977 7228 4983
rect 7364 4977 7900 4983
rect 7924 4977 7948 4983
rect 36 4957 188 4963
rect 260 4957 316 4963
rect 324 4957 428 4963
rect 468 4957 556 4963
rect 564 4957 828 4963
rect 1012 4957 1196 4963
rect 1204 4957 1420 4963
rect 1428 4957 1580 4963
rect 2132 4957 2220 4963
rect 2228 4957 2492 4963
rect 2500 4957 2668 4963
rect 2676 4957 3004 4963
rect 3236 4957 3324 4963
rect 3348 4957 3388 4963
rect 3396 4957 3420 4963
rect 3444 4957 4124 4963
rect 4164 4957 4716 4963
rect 6036 4957 7036 4963
rect 7620 4957 7788 4963
rect 7796 4957 7932 4963
rect 7940 4957 7996 4963
rect 20 4937 44 4943
rect 52 4937 268 4943
rect 276 4937 284 4943
rect 372 4937 412 4943
rect 820 4937 860 4943
rect 868 4937 1612 4943
rect 1620 4937 1804 4943
rect 1812 4937 1820 4943
rect 1940 4937 1964 4943
rect 2356 4937 2364 4943
rect 2372 4937 2396 4943
rect 2404 4937 2428 4943
rect 2436 4937 2444 4943
rect 2452 4937 2540 4943
rect 2548 4937 2636 4943
rect 2644 4937 2684 4943
rect 2740 4937 2796 4943
rect 2820 4937 2892 4943
rect 3028 4937 3500 4943
rect 3508 4937 3580 4943
rect 3588 4937 3612 4943
rect 4596 4937 4764 4943
rect 4980 4937 5068 4943
rect 5412 4937 5564 4943
rect 5652 4937 5740 4943
rect 5972 4937 6060 4943
rect 6116 4937 6300 4943
rect 6788 4937 6860 4943
rect 6932 4937 7036 4943
rect 7268 4937 7516 4943
rect 7684 4937 7740 4943
rect 7748 4937 7932 4943
rect 8004 4937 8092 4943
rect 84 4917 268 4923
rect 292 4917 460 4923
rect 612 4917 636 4923
rect 884 4917 1148 4923
rect 1204 4917 1260 4923
rect 1316 4917 1452 4923
rect 1508 4917 1580 4923
rect 2244 4917 2300 4923
rect 2452 4917 2524 4923
rect 2580 4917 2636 4923
rect 2708 4917 3148 4923
rect 3380 4917 3564 4923
rect 3572 4917 3676 4923
rect 3876 4917 3980 4923
rect 4260 4917 4364 4923
rect 5204 4917 5212 4923
rect 5460 4917 5676 4923
rect 5700 4917 5756 4923
rect 5764 4917 6220 4923
rect 6436 4917 6492 4923
rect 6676 4917 6700 4923
rect 6804 4917 6924 4923
rect 6980 4917 7116 4923
rect 7236 4917 7244 4923
rect 7556 4917 7660 4923
rect 7732 4917 7772 4923
rect 180 4897 220 4903
rect 260 4897 348 4903
rect 404 4897 460 4903
rect 564 4897 604 4903
rect 644 4897 716 4903
rect 1236 4897 1436 4903
rect 1444 4897 1516 4903
rect 2100 4897 2140 4903
rect 2180 4897 2220 4903
rect 2228 4897 2300 4903
rect 2340 4897 2380 4903
rect 2573 4903 2579 4916
rect 2388 4897 2579 4903
rect 2660 4897 2764 4903
rect 2788 4897 2828 4903
rect 2868 4897 2972 4903
rect 3172 4897 3180 4903
rect 3556 4897 3884 4903
rect 4372 4897 4620 4903
rect 5364 4897 5436 4903
rect 5732 4897 5756 4903
rect 6436 4897 6652 4903
rect 6701 4903 6707 4916
rect 6701 4897 6876 4903
rect 6884 4897 6908 4903
rect 6916 4897 6956 4903
rect 7652 4897 7692 4903
rect 7780 4897 7868 4903
rect 100 4877 156 4883
rect 164 4877 380 4883
rect 436 4877 508 4883
rect 532 4877 572 4883
rect 580 4877 588 4883
rect 660 4877 892 4883
rect 1332 4877 1596 4883
rect 2020 4877 2140 4883
rect 2180 4877 2252 4883
rect 2404 4877 2460 4883
rect 2532 4877 2876 4883
rect 3220 4877 3228 4883
rect 3428 4877 3484 4883
rect 3492 4877 3532 4883
rect 3716 4877 3804 4883
rect 3828 4877 4140 4883
rect 4724 4877 4748 4883
rect 4756 4877 4796 4883
rect 5140 4877 5452 4883
rect 5556 4877 5788 4883
rect 6628 4877 6668 4883
rect 6756 4877 6892 4883
rect 6932 4877 7084 4883
rect 7620 4877 7836 4883
rect 7972 4877 8044 4883
rect 8052 4877 8124 4883
rect 564 4857 748 4863
rect 756 4857 844 4863
rect 1364 4857 1468 4863
rect 2164 4857 2380 4863
rect 3156 4857 3356 4863
rect 3412 4857 3468 4863
rect 3476 4857 3676 4863
rect 5476 4857 5548 4863
rect 5588 4857 5820 4863
rect 6164 4857 6220 4863
rect 7652 4857 7724 4863
rect 7908 4857 8108 4863
rect 308 4837 412 4843
rect 420 4837 700 4843
rect 1732 4837 1980 4843
rect 3204 4837 4156 4843
rect 4164 4837 4396 4843
rect 4404 4837 4604 4843
rect 5012 4837 5052 4843
rect 5252 4837 5404 4843
rect 5716 4837 6204 4843
rect 6324 4837 6572 4843
rect 7636 4837 7692 4843
rect 452 4817 620 4823
rect 3956 4817 4108 4823
rect 4116 4817 4444 4823
rect 4948 4817 5148 4823
rect 1736 4814 1784 4816
rect 1736 4806 1740 4814
rect 1750 4806 1756 4814
rect 1764 4806 1770 4814
rect 1780 4806 1784 4814
rect 1736 4804 1784 4806
rect 4808 4814 4856 4816
rect 4808 4806 4812 4814
rect 4822 4806 4828 4814
rect 4836 4806 4842 4814
rect 4852 4806 4856 4814
rect 4808 4804 4856 4806
rect 1460 4797 1484 4803
rect 2100 4797 2572 4803
rect 2580 4797 2668 4803
rect 3172 4797 3836 4803
rect 4356 4797 4636 4803
rect 7876 4797 7964 4803
rect 180 4777 524 4783
rect 532 4777 684 4783
rect 692 4777 716 4783
rect 1204 4777 1292 4783
rect 1300 4777 1644 4783
rect 2244 4777 3132 4783
rect 3556 4777 3708 4783
rect 4292 4777 4476 4783
rect 4500 4777 6028 4783
rect 7284 4777 7596 4783
rect 292 4757 764 4763
rect 1316 4757 1628 4763
rect 2468 4757 2860 4763
rect 3629 4757 3820 4763
rect 3629 4744 3635 4757
rect 4452 4757 4476 4763
rect 4916 4757 5004 4763
rect 5028 4757 5052 4763
rect 5124 4757 5164 4763
rect 5444 4757 5516 4763
rect 6052 4757 6684 4763
rect 6692 4757 6732 4763
rect 6740 4757 6828 4763
rect 6900 4757 7068 4763
rect 7524 4757 7708 4763
rect 7716 4757 7852 4763
rect 7972 4757 8092 4763
rect 196 4737 300 4743
rect 372 4737 460 4743
rect 676 4737 812 4743
rect 1444 4737 1820 4743
rect 2052 4737 2124 4743
rect 2292 4737 2588 4743
rect 2740 4737 2828 4743
rect 3604 4737 3628 4743
rect 3732 4737 3772 4743
rect 4116 4737 6076 4743
rect 6084 4737 6460 4743
rect 6468 4737 6844 4743
rect 6852 4737 6876 4743
rect 6884 4737 6908 4743
rect 7540 4737 7676 4743
rect 7684 4737 7756 4743
rect 7764 4737 7884 4743
rect 276 4717 348 4723
rect 356 4717 476 4723
rect 660 4717 684 4723
rect 836 4717 876 4723
rect 980 4717 1132 4723
rect 1268 4717 1388 4723
rect 1492 4717 1820 4723
rect 2116 4717 2412 4723
rect 2596 4717 2796 4723
rect 2852 4717 3052 4723
rect 3124 4717 3196 4723
rect 3604 4717 3692 4723
rect 3940 4717 3996 4723
rect 4004 4717 4156 4723
rect 4740 4717 4828 4723
rect 4836 4717 4940 4723
rect 4948 4717 4988 4723
rect 4996 4717 5036 4723
rect 5060 4717 5180 4723
rect 5284 4717 5340 4723
rect 5364 4717 5388 4723
rect 5460 4717 5532 4723
rect 5540 4717 5932 4723
rect 5940 4717 5964 4723
rect 6212 4717 6236 4723
rect 6564 4717 6652 4723
rect 6660 4717 6732 4723
rect 6740 4717 6812 4723
rect 6868 4717 6956 4723
rect 7300 4717 7436 4723
rect 7588 4717 7692 4723
rect 7700 4717 7820 4723
rect 8004 4717 8060 4723
rect 148 4697 268 4703
rect 372 4697 396 4703
rect 404 4697 588 4703
rect 596 4697 636 4703
rect 644 4697 732 4703
rect 740 4697 1852 4703
rect 2132 4697 2172 4703
rect 2372 4697 2444 4703
rect 2484 4697 2524 4703
rect 2772 4697 2924 4703
rect 2932 4697 3356 4703
rect 3428 4697 3516 4703
rect 3572 4697 3868 4703
rect 3988 4697 4012 4703
rect 4356 4697 4492 4703
rect 4564 4697 4588 4703
rect 4612 4697 4684 4703
rect 4708 4697 4716 4703
rect 4724 4697 4748 4703
rect 4756 4697 5100 4703
rect 5332 4697 5340 4703
rect 5476 4697 5500 4703
rect 5524 4697 5596 4703
rect 5636 4697 5676 4703
rect 5684 4697 5852 4703
rect 5860 4697 5932 4703
rect 6020 4697 6156 4703
rect 6164 4697 6316 4703
rect 6324 4697 6700 4703
rect 6708 4697 6748 4703
rect 6804 4697 6924 4703
rect 6964 4697 7036 4703
rect 7412 4697 7484 4703
rect 7492 4697 7548 4703
rect 7668 4697 7692 4703
rect 7700 4697 7804 4703
rect 7860 4697 7948 4703
rect 7956 4697 8012 4703
rect 228 4677 572 4683
rect 580 4677 652 4683
rect 724 4677 940 4683
rect 1188 4677 1292 4683
rect 1300 4677 1452 4683
rect 1460 4677 1500 4683
rect 1588 4677 1628 4683
rect 1636 4677 1900 4683
rect 2084 4677 2108 4683
rect 2228 4677 2460 4683
rect 2804 4677 2972 4683
rect 3188 4677 3228 4683
rect 3236 4677 3404 4683
rect 3572 4677 3644 4683
rect 3652 4677 3772 4683
rect 4221 4683 4227 4696
rect 3972 4677 4227 4683
rect 4372 4677 4412 4683
rect 4420 4677 4460 4683
rect 4468 4677 4524 4683
rect 4564 4677 4684 4683
rect 4692 4677 4764 4683
rect 4772 4677 5116 4683
rect 5124 4677 5164 4683
rect 5220 4677 5644 4683
rect 5652 4677 5724 4683
rect 5748 4677 5820 4683
rect 6164 4677 6220 4683
rect 6228 4677 6284 4683
rect 6420 4677 6604 4683
rect 6612 4677 6636 4683
rect 6820 4677 7084 4683
rect 7092 4677 7132 4683
rect 7140 4677 7180 4683
rect 7572 4677 7612 4683
rect 7828 4677 7884 4683
rect 7892 4677 7916 4683
rect 260 4657 316 4663
rect 1140 4657 1260 4663
rect 1332 4657 1388 4663
rect 1540 4657 1708 4663
rect 2164 4657 2252 4663
rect 2436 4657 2492 4663
rect 3076 4657 3164 4663
rect 3540 4657 3580 4663
rect 3684 4657 3756 4663
rect 4365 4663 4371 4676
rect 3908 4657 4371 4663
rect 4516 4657 4572 4663
rect 4596 4657 4652 4663
rect 4676 4657 4748 4663
rect 4756 4657 4860 4663
rect 4868 4657 4972 4663
rect 4980 4657 5036 4663
rect 5332 4657 5452 4663
rect 5492 4657 5548 4663
rect 5556 4657 5708 4663
rect 5716 4657 5788 4663
rect 5956 4657 6396 4663
rect 6404 4657 6476 4663
rect 6516 4657 6540 4663
rect 6580 4657 6796 4663
rect 6996 4657 7100 4663
rect 7156 4657 7164 4663
rect 7636 4657 7676 4663
rect 7684 4657 7740 4663
rect 7796 4657 7852 4663
rect 7924 4657 8028 4663
rect 8068 4657 8083 4663
rect 8077 4644 8083 4657
rect 20 4637 60 4643
rect 68 4637 204 4643
rect 260 4637 284 4643
rect 292 4637 604 4643
rect 628 4637 1116 4643
rect 1124 4637 2044 4643
rect 2100 4637 2140 4643
rect 2148 4637 2300 4643
rect 2308 4637 2380 4643
rect 2388 4637 2588 4643
rect 2596 4637 3276 4643
rect 3924 4637 4060 4643
rect 4068 4637 4348 4643
rect 4452 4637 4636 4643
rect 5204 4637 5260 4643
rect 5348 4637 5692 4643
rect 5700 4637 5756 4643
rect 6116 4637 6140 4643
rect 6180 4637 6364 4643
rect 6532 4637 6620 4643
rect 7732 4637 7788 4643
rect 868 4617 908 4623
rect 916 4617 3244 4623
rect 3700 4617 3948 4623
rect 4100 4617 4412 4623
rect 4452 4617 4764 4623
rect 5060 4617 5500 4623
rect 5508 4617 5772 4623
rect 5780 4617 5884 4623
rect 7572 4617 7692 4623
rect 7716 4617 7900 4623
rect 8052 4617 8124 4623
rect 3272 4614 3320 4616
rect 3272 4606 3276 4614
rect 3286 4606 3292 4614
rect 3300 4606 3306 4614
rect 3316 4606 3320 4614
rect 3272 4604 3320 4606
rect 6344 4614 6392 4616
rect 6344 4606 6348 4614
rect 6358 4606 6364 4614
rect 6372 4606 6378 4614
rect 6388 4606 6392 4614
rect 6344 4604 6392 4606
rect 868 4597 972 4603
rect 1332 4597 1420 4603
rect 1428 4597 1468 4603
rect 1476 4597 1548 4603
rect 1828 4597 1916 4603
rect 1924 4597 2060 4603
rect 2484 4597 2812 4603
rect 3732 4597 3916 4603
rect 4244 4597 4380 4603
rect 4580 4597 4588 4603
rect 5277 4597 5731 4603
rect 324 4577 348 4583
rect 788 4577 812 4583
rect 1012 4577 1100 4583
rect 1812 4577 1852 4583
rect 1860 4577 3228 4583
rect 3252 4577 3292 4583
rect 3876 4577 3900 4583
rect 3908 4577 3948 4583
rect 3956 4577 4044 4583
rect 4052 4577 4220 4583
rect 4340 4577 4428 4583
rect 5277 4583 5283 4597
rect 4516 4577 5283 4583
rect 5508 4577 5628 4583
rect 5668 4577 5692 4583
rect 5725 4583 5731 4597
rect 5780 4597 5868 4603
rect 5940 4597 5996 4603
rect 7556 4597 7580 4603
rect 8004 4597 8028 4603
rect 5725 4577 5948 4583
rect 6452 4577 6492 4583
rect 6500 4577 6620 4583
rect 6628 4577 6796 4583
rect 7444 4577 7564 4583
rect 308 4557 524 4563
rect 1540 4557 1596 4563
rect 1620 4557 1740 4563
rect 2420 4557 2540 4563
rect 2548 4557 2684 4563
rect 2708 4557 2764 4563
rect 2836 4557 2860 4563
rect 3332 4557 3564 4563
rect 3652 4557 3852 4563
rect 4509 4563 4515 4576
rect 4324 4557 4515 4563
rect 5092 4557 5228 4563
rect 5684 4557 5756 4563
rect 5892 4557 6092 4563
rect 6292 4557 6492 4563
rect 6532 4557 6636 4563
rect 6708 4557 6828 4563
rect 7204 4557 7276 4563
rect 7364 4557 7404 4563
rect 7412 4557 7484 4563
rect 7556 4557 7580 4563
rect 7732 4557 7772 4563
rect 420 4537 476 4543
rect 1588 4537 1692 4543
rect 2148 4537 2364 4543
rect 2372 4537 2396 4543
rect 2404 4537 2716 4543
rect 2724 4537 2876 4543
rect 2980 4537 3084 4543
rect 3156 4537 3180 4543
rect 3220 4537 3244 4543
rect 3780 4537 3852 4543
rect 3924 4537 4028 4543
rect 4036 4537 4092 4543
rect 4260 4537 4284 4543
rect 4292 4537 4348 4543
rect 5076 4537 5116 4543
rect 5124 4537 5180 4543
rect 5396 4537 5548 4543
rect 5620 4537 5660 4543
rect 5732 4537 5884 4543
rect 6052 4537 6252 4543
rect 6612 4537 6764 4543
rect 6788 4537 6828 4543
rect 6836 4537 6908 4543
rect 7172 4537 7372 4543
rect 7476 4537 7532 4543
rect 7540 4537 7612 4543
rect 7716 4537 7852 4543
rect 7924 4537 8012 4543
rect 244 4517 364 4523
rect 372 4517 444 4523
rect 516 4517 684 4523
rect 836 4517 988 4523
rect 1076 4517 1132 4523
rect 1588 4517 1676 4523
rect 1748 4517 1820 4523
rect 1828 4517 1980 4523
rect 1988 4517 2204 4523
rect 2276 4517 2332 4523
rect 2452 4517 2492 4523
rect 2532 4517 2748 4523
rect 2756 4517 2860 4523
rect 2973 4523 2979 4536
rect 2868 4517 2979 4523
rect 3588 4517 3612 4523
rect 3668 4517 3948 4523
rect 4004 4517 4028 4523
rect 4180 4517 4268 4523
rect 4324 4517 4348 4523
rect 4612 4517 4620 4523
rect 4628 4517 4684 4523
rect 4692 4517 4924 4523
rect 4932 4517 5132 4523
rect 5540 4517 5564 4523
rect 5636 4517 5756 4523
rect 5828 4517 5884 4523
rect 6228 4517 6540 4523
rect 6692 4517 6972 4523
rect 7172 4517 7228 4523
rect 7652 4517 7740 4523
rect 7748 4517 7836 4523
rect 7988 4517 8060 4523
rect 308 4497 380 4503
rect 420 4497 684 4503
rect 900 4497 1020 4503
rect 1028 4497 1164 4503
rect 1508 4497 1612 4503
rect 2132 4497 2140 4503
rect 2372 4497 2460 4503
rect 2493 4503 2499 4516
rect 2493 4497 2540 4503
rect 2692 4497 2716 4503
rect 2804 4497 2908 4503
rect 2932 4497 3036 4503
rect 3412 4497 3676 4503
rect 3796 4497 3804 4503
rect 3812 4497 3980 4503
rect 3988 4497 4188 4503
rect 4564 4497 5052 4503
rect 5412 4497 5580 4503
rect 5588 4497 5724 4503
rect 6212 4497 6284 4503
rect 6420 4497 6556 4503
rect 6660 4497 6844 4503
rect 6852 4497 6860 4503
rect 7284 4497 7372 4503
rect 452 4477 508 4483
rect 1060 4477 1084 4483
rect 1604 4477 2220 4483
rect 2356 4477 2412 4483
rect 2452 4477 2540 4483
rect 2676 4477 2796 4483
rect 3236 4477 3436 4483
rect 3524 4477 3820 4483
rect 4564 4477 4780 4483
rect 4980 4477 5068 4483
rect 5332 4477 5516 4483
rect 5572 4477 5612 4483
rect 6068 4477 6108 4483
rect 6532 4477 6668 4483
rect 6756 4477 7100 4483
rect 7108 4477 7292 4483
rect 7940 4477 8124 4483
rect 1044 4457 1132 4463
rect 2004 4457 2044 4463
rect 2669 4463 2675 4476
rect 2388 4457 2675 4463
rect 3821 4463 3827 4476
rect 3821 4457 3964 4463
rect 3972 4457 4012 4463
rect 4020 4457 4108 4463
rect 4724 4457 4876 4463
rect 5188 4457 6124 4463
rect 6132 4457 6140 4463
rect 1348 4437 1388 4443
rect 2052 4437 2108 4443
rect 3172 4437 3196 4443
rect 3204 4437 3260 4443
rect 3268 4437 3868 4443
rect 3972 4437 4076 4443
rect 4148 4437 4460 4443
rect 4644 4437 4732 4443
rect 4740 4437 4844 4443
rect 4852 4437 4876 4443
rect 5012 4437 5420 4443
rect 5956 4437 6748 4443
rect 7060 4437 7132 4443
rect 7156 4437 7484 4443
rect 8004 4437 8092 4443
rect 3364 4417 4300 4423
rect 4996 4417 5052 4423
rect 5300 4417 5804 4423
rect 7156 4417 7196 4423
rect 7428 4417 7532 4423
rect 1736 4414 1784 4416
rect 1736 4406 1740 4414
rect 1750 4406 1756 4414
rect 1764 4406 1770 4414
rect 1780 4406 1784 4414
rect 1736 4404 1784 4406
rect 4808 4414 4856 4416
rect 4808 4406 4812 4414
rect 4822 4406 4828 4414
rect 4836 4406 4842 4414
rect 4852 4406 4856 4414
rect 4808 4404 4856 4406
rect 20 4397 108 4403
rect 932 4397 956 4403
rect 2436 4397 3164 4403
rect 4052 4397 4076 4403
rect 5236 4397 5836 4403
rect 7460 4397 7516 4403
rect 7588 4397 7948 4403
rect 7956 4397 8060 4403
rect 2884 4377 4044 4383
rect 148 4357 300 4363
rect 356 4357 780 4363
rect 996 4357 1148 4363
rect 1156 4357 1260 4363
rect 1268 4357 1356 4363
rect 2820 4357 3004 4363
rect 3956 4357 4220 4363
rect 5588 4357 5756 4363
rect 5764 4357 5884 4363
rect 6029 4357 6300 4363
rect 6029 4344 6035 4357
rect 7444 4357 7564 4363
rect 7636 4357 7900 4363
rect 244 4337 700 4343
rect 2084 4337 2204 4343
rect 2244 4337 2268 4343
rect 2708 4337 2908 4343
rect 3844 4337 3868 4343
rect 3892 4337 4012 4343
rect 4020 4337 4060 4343
rect 4324 4337 4460 4343
rect 4484 4337 5132 4343
rect 5140 4337 5180 4343
rect 5476 4337 5708 4343
rect 5748 4337 5868 4343
rect 5972 4337 6028 4343
rect 6084 4337 6124 4343
rect 6164 4337 6355 4343
rect 6349 4324 6355 4337
rect 6692 4337 6748 4343
rect 6804 4337 6956 4343
rect 7124 4337 7196 4343
rect 7204 4337 7292 4343
rect 7300 4337 7500 4343
rect 7700 4337 7756 4343
rect 7780 4337 7804 4343
rect 180 4317 284 4323
rect 308 4317 428 4323
rect 596 4317 636 4323
rect 692 4317 732 4323
rect 1028 4317 1052 4323
rect 1412 4317 1500 4323
rect 1668 4317 1916 4323
rect 2100 4317 2156 4323
rect 2164 4317 2396 4323
rect 2884 4317 2940 4323
rect 3428 4317 3996 4323
rect 4004 4317 4284 4323
rect 4292 4317 4444 4323
rect 4580 4317 4588 4323
rect 4900 4317 5532 4323
rect 5789 4317 6204 4323
rect 5789 4304 5795 4317
rect 6212 4317 6236 4323
rect 6292 4317 6316 4323
rect 6356 4317 6524 4323
rect 6701 4317 6860 4323
rect 6701 4304 6707 4317
rect 7124 4317 7244 4323
rect 7268 4317 7324 4323
rect 7364 4317 7388 4323
rect 7444 4317 7596 4323
rect 7684 4317 7740 4323
rect 7748 4317 7820 4323
rect 228 4297 348 4303
rect 484 4297 524 4303
rect 580 4297 828 4303
rect 980 4297 1100 4303
rect 1108 4297 1228 4303
rect 1236 4297 1292 4303
rect 1444 4297 1548 4303
rect 1716 4297 1772 4303
rect 1844 4297 2316 4303
rect 2468 4297 2556 4303
rect 2788 4297 2844 4303
rect 2996 4297 3020 4303
rect 3460 4297 3484 4303
rect 3540 4297 3612 4303
rect 4084 4297 4188 4303
rect 4596 4297 4652 4303
rect 4708 4297 4844 4303
rect 4996 4297 5260 4303
rect 5268 4297 5308 4303
rect 5572 4297 5612 4303
rect 5620 4297 5660 4303
rect 5732 4297 5788 4303
rect 6084 4297 6380 4303
rect 6612 4297 6700 4303
rect 6852 4297 6908 4303
rect 7204 4297 7276 4303
rect 7380 4297 7452 4303
rect 7556 4297 7628 4303
rect 7780 4297 7836 4303
rect 8004 4297 8028 4303
rect 164 4277 236 4283
rect 388 4277 412 4283
rect 420 4277 636 4283
rect 644 4277 732 4283
rect 740 4277 780 4283
rect 788 4277 828 4283
rect 1060 4277 1132 4283
rect 1140 4277 1180 4283
rect 1204 4277 1244 4283
rect 1444 4277 1452 4283
rect 1540 4277 1612 4283
rect 2004 4277 2076 4283
rect 2500 4277 2716 4283
rect 2724 4277 2764 4283
rect 2772 4277 2812 4283
rect 2941 4277 3068 4283
rect 36 4257 236 4263
rect 516 4257 636 4263
rect 820 4257 860 4263
rect 1044 4257 1116 4263
rect 1124 4257 1292 4263
rect 1300 4257 1324 4263
rect 1332 4257 1404 4263
rect 1540 4257 1628 4263
rect 1716 4257 1868 4263
rect 2148 4257 2252 4263
rect 2404 4257 2460 4263
rect 2941 4263 2947 4277
rect 3140 4277 3436 4283
rect 3540 4277 3628 4283
rect 3796 4277 3948 4283
rect 4324 4277 4988 4283
rect 5044 4277 5052 4283
rect 5060 4277 5148 4283
rect 5556 4277 5708 4283
rect 5764 4277 5804 4283
rect 5876 4277 5980 4283
rect 5988 4277 6172 4283
rect 6308 4277 6444 4283
rect 6692 4277 6716 4283
rect 6836 4277 6892 4283
rect 7236 4277 7260 4283
rect 7316 4277 7468 4283
rect 7780 4277 7820 4283
rect 2692 4257 2947 4263
rect 3028 4257 3052 4263
rect 3060 4257 3260 4263
rect 3268 4257 3324 4263
rect 3444 4257 4508 4263
rect 4532 4257 4972 4263
rect 5028 4257 5212 4263
rect 5220 4257 5244 4263
rect 5796 4257 5900 4263
rect 5908 4257 5996 4263
rect 6148 4257 6204 4263
rect 6324 4257 6412 4263
rect 6500 4257 6588 4263
rect 7124 4257 7212 4263
rect 7236 4257 7436 4263
rect 7460 4257 7580 4263
rect 7684 4257 7964 4263
rect 36 4237 252 4243
rect 493 4243 499 4256
rect 493 4237 540 4243
rect 1876 4237 1964 4243
rect 1972 4237 2156 4243
rect 2164 4237 2204 4243
rect 2724 4237 2828 4243
rect 3028 4237 3148 4243
rect 3172 4237 3292 4243
rect 3620 4237 3724 4243
rect 3732 4237 3756 4243
rect 3764 4237 3804 4243
rect 3876 4237 3948 4243
rect 3956 4237 4700 4243
rect 4740 4237 4780 4243
rect 4868 4237 4956 4243
rect 4964 4237 5052 4243
rect 5204 4237 5404 4243
rect 5412 4237 5596 4243
rect 5652 4237 5836 4243
rect 5997 4243 6003 4256
rect 5997 4237 6188 4243
rect 6436 4237 6620 4243
rect 7140 4237 7148 4243
rect 7213 4243 7219 4256
rect 7213 4237 7388 4243
rect 7396 4237 7500 4243
rect 116 4217 252 4223
rect 260 4217 332 4223
rect 340 4217 508 4223
rect 1988 4217 2412 4223
rect 2596 4217 2924 4223
rect 3060 4217 3116 4223
rect 3805 4223 3811 4236
rect 3805 4217 4124 4223
rect 4733 4223 4739 4236
rect 4516 4217 4739 4223
rect 4772 4217 4940 4223
rect 5092 4217 5244 4223
rect 5604 4217 5820 4223
rect 5876 4217 5932 4223
rect 6148 4217 6252 4223
rect 6564 4217 6652 4223
rect 6788 4217 6924 4223
rect 7092 4217 7260 4223
rect 7268 4217 7372 4223
rect 7716 4217 7788 4223
rect 3272 4214 3320 4216
rect 3272 4206 3276 4214
rect 3286 4206 3292 4214
rect 3300 4206 3306 4214
rect 3316 4206 3320 4214
rect 3272 4204 3320 4206
rect 6344 4214 6392 4216
rect 6344 4206 6348 4214
rect 6358 4206 6364 4214
rect 6372 4206 6378 4214
rect 6388 4206 6392 4214
rect 6344 4204 6392 4206
rect 196 4197 204 4203
rect 276 4197 364 4203
rect 1140 4197 1388 4203
rect 2116 4197 2428 4203
rect 2548 4197 2700 4203
rect 2884 4197 2924 4203
rect 3012 4197 3212 4203
rect 3572 4197 4012 4203
rect 4020 4197 4188 4203
rect 4276 4197 4396 4203
rect 4404 4197 4492 4203
rect 4516 4197 4844 4203
rect 5012 4197 5068 4203
rect 5124 4197 5324 4203
rect 5332 4197 5452 4203
rect 5860 4197 6204 4203
rect 6468 4197 6492 4203
rect 6580 4197 6652 4203
rect 6669 4197 6972 4203
rect 436 4177 492 4183
rect 836 4177 876 4183
rect 1012 4177 1436 4183
rect 1725 4177 1836 4183
rect 1725 4164 1731 4177
rect 1844 4177 1852 4183
rect 1908 4177 3180 4183
rect 3396 4177 3772 4183
rect 3796 4177 4028 4183
rect 4452 4177 4556 4183
rect 4564 4177 4860 4183
rect 4932 4177 4972 4183
rect 5188 4177 5228 4183
rect 5284 4177 5468 4183
rect 5764 4177 5852 4183
rect 5860 4177 6076 4183
rect 6148 4177 6188 4183
rect 6196 4177 6492 4183
rect 6669 4183 6675 4197
rect 7380 4197 7564 4203
rect 8036 4197 8076 4203
rect 6532 4177 6675 4183
rect 7108 4177 7308 4183
rect 7764 4177 7948 4183
rect 8052 4177 8060 4183
rect 180 4157 204 4163
rect 916 4157 1052 4163
rect 1252 4157 1452 4163
rect 1460 4157 1516 4163
rect 1588 4157 1724 4163
rect 1764 4157 1916 4163
rect 1924 4157 2012 4163
rect 2020 4157 2268 4163
rect 2628 4157 2684 4163
rect 2916 4157 2988 4163
rect 3364 4157 3644 4163
rect 3652 4157 3708 4163
rect 3764 4157 3916 4163
rect 4164 4157 4348 4163
rect 4388 4157 4412 4163
rect 4548 4157 4716 4163
rect 4724 4157 4796 4163
rect 4948 4157 5340 4163
rect 5524 4157 5692 4163
rect 5700 4157 5740 4163
rect 5764 4157 5820 4163
rect 6020 4157 6268 4163
rect 6324 4157 6668 4163
rect 6692 4157 6844 4163
rect 7316 4157 7388 4163
rect 7444 4157 7468 4163
rect 7652 4157 7708 4163
rect 7844 4157 7900 4163
rect 8052 4157 8124 4163
rect 8132 4157 8140 4163
rect 148 4137 188 4143
rect 484 4137 716 4143
rect 900 4137 940 4143
rect 948 4137 956 4143
rect 964 4137 1100 4143
rect 1108 4137 1436 4143
rect 1444 4137 1500 4143
rect 1508 4137 1596 4143
rect 1604 4137 1820 4143
rect 1828 4137 1932 4143
rect 1940 4137 2028 4143
rect 2036 4137 2140 4143
rect 2324 4137 2476 4143
rect 3188 4137 3340 4143
rect 3348 4137 3372 4143
rect 3476 4137 3500 4143
rect 3780 4137 4684 4143
rect 4708 4137 4780 4143
rect 4884 4137 4892 4143
rect 4980 4137 5356 4143
rect 5364 4137 5372 4143
rect 5652 4137 5868 4143
rect 6052 4137 6252 4143
rect 6484 4137 6684 4143
rect 6996 4137 7100 4143
rect 7188 4137 7228 4143
rect 7284 4137 7324 4143
rect 7332 4137 7372 4143
rect 7524 4137 7708 4143
rect 7716 4137 8012 4143
rect 8020 4137 8076 4143
rect 196 4117 284 4123
rect 692 4117 748 4123
rect 1044 4117 1116 4123
rect 1172 4117 1356 4123
rect 1380 4117 1436 4123
rect 1508 4117 1612 4123
rect 1636 4117 2044 4123
rect 2052 4117 2188 4123
rect 2244 4117 2444 4123
rect 2516 4117 2588 4123
rect 2596 4117 2636 4123
rect 2676 4117 2716 4123
rect 2788 4117 2812 4123
rect 2836 4117 2956 4123
rect 3332 4117 3484 4123
rect 3684 4117 3724 4123
rect 3732 4117 3772 4123
rect 3828 4117 3948 4123
rect 4020 4117 4300 4123
rect 4308 4117 4332 4123
rect 4372 4117 4492 4123
rect 4548 4117 4988 4123
rect 5044 4117 5116 4123
rect 5181 4117 5276 4123
rect 68 4097 140 4103
rect 596 4097 636 4103
rect 1012 4097 1068 4103
rect 1124 4097 1148 4103
rect 1572 4097 1644 4103
rect 1908 4097 1932 4103
rect 2196 4097 2364 4103
rect 2708 4097 2764 4103
rect 2804 4097 2908 4103
rect 2980 4097 3084 4103
rect 3204 4097 3532 4103
rect 3924 4097 3996 4103
rect 4244 4097 5020 4103
rect 5181 4103 5187 4117
rect 5300 4117 5356 4123
rect 5396 4117 5420 4123
rect 5620 4117 5772 4123
rect 5780 4117 6076 4123
rect 6084 4117 6300 4123
rect 6516 4117 6748 4123
rect 6756 4117 6812 4123
rect 7108 4117 7196 4123
rect 7252 4117 7308 4123
rect 7332 4117 7356 4123
rect 7556 4117 7900 4123
rect 8116 4117 8140 4123
rect 5108 4097 5187 4103
rect 5204 4097 5308 4103
rect 5572 4097 5660 4103
rect 5700 4097 5724 4103
rect 6628 4097 6668 4103
rect 6708 4097 6748 4103
rect 7188 4097 7404 4103
rect 7620 4097 7660 4103
rect 7668 4097 8092 4103
rect 1092 4077 1164 4083
rect 1428 4077 2844 4083
rect 2884 4077 2940 4083
rect 3492 4077 3884 4083
rect 3892 4077 4460 4083
rect 4468 4077 4508 4083
rect 4516 4077 4588 4083
rect 4596 4077 4748 4083
rect 5044 4077 5068 4083
rect 5092 4077 6972 4083
rect 6980 4077 7164 4083
rect 7172 4077 7452 4083
rect 7460 4077 7468 4083
rect 7748 4077 7788 4083
rect 7796 4077 7804 4083
rect 7972 4077 8012 4083
rect 548 4057 1148 4063
rect 1540 4057 1996 4063
rect 2004 4057 2316 4063
rect 2500 4057 2684 4063
rect 2692 4057 3692 4063
rect 4084 4057 4316 4063
rect 4692 4057 4876 4063
rect 4900 4057 5180 4063
rect 5380 4057 5820 4063
rect 6724 4057 6844 4063
rect 7748 4057 7804 4063
rect 7821 4057 7868 4063
rect 692 4037 732 4043
rect 932 4037 1020 4043
rect 1028 4037 1084 4043
rect 1092 4037 1260 4043
rect 1892 4037 3676 4043
rect 3693 4043 3699 4056
rect 3693 4037 5916 4043
rect 5924 4037 6204 4043
rect 6212 4037 6828 4043
rect 7620 4037 7772 4043
rect 7821 4043 7827 4057
rect 7908 4057 7964 4063
rect 7812 4037 7827 4043
rect 7844 4037 8044 4043
rect 84 4017 316 4023
rect 324 4017 444 4023
rect 452 4017 476 4023
rect 2340 4017 2380 4023
rect 2532 4017 2604 4023
rect 2612 4017 2780 4023
rect 2852 4017 3324 4023
rect 3540 4017 3932 4023
rect 3988 4017 4540 4023
rect 4884 4017 5052 4023
rect 5060 4017 5212 4023
rect 5236 4017 5628 4023
rect 5828 4017 7180 4023
rect 7828 4017 8092 4023
rect 1736 4014 1784 4016
rect 1736 4006 1740 4014
rect 1750 4006 1756 4014
rect 1764 4006 1770 4014
rect 1780 4006 1784 4014
rect 1736 4004 1784 4006
rect 4808 4014 4856 4016
rect 4808 4006 4812 4014
rect 4822 4006 4828 4014
rect 4836 4006 4842 4014
rect 4852 4006 4856 4014
rect 4808 4004 4856 4006
rect 2276 3997 2636 4003
rect 2724 3997 2764 4003
rect 2772 3997 2988 4003
rect 3396 3997 3468 4003
rect 3668 3997 3772 4003
rect 4068 3997 4268 4003
rect 4324 3997 4348 4003
rect 4484 3997 4668 4003
rect 4676 3997 4748 4003
rect 5236 3997 5276 4003
rect 5508 3997 5612 4003
rect 5668 3997 5884 4003
rect 5892 3997 6108 4003
rect 6356 3997 6668 4003
rect 7892 3997 8092 4003
rect 868 3977 1324 3983
rect 1332 3977 1420 3983
rect 2452 3977 3132 3983
rect 3412 3977 3484 3983
rect 3508 3977 3548 3983
rect 3556 3977 4028 3983
rect 4036 3977 4412 3983
rect 4420 3977 6428 3983
rect 7316 3977 7596 3983
rect 7892 3977 7996 3983
rect 548 3957 940 3963
rect 2548 3957 2572 3963
rect 2580 3957 2700 3963
rect 3220 3957 4364 3963
rect 4372 3957 4732 3963
rect 5460 3957 6268 3963
rect 6276 3957 6540 3963
rect 6740 3957 7612 3963
rect 7748 3957 7788 3963
rect 7796 3957 7980 3963
rect 7988 3957 7996 3963
rect 8004 3957 8108 3963
rect 292 3937 572 3943
rect 580 3937 1100 3943
rect 1700 3937 1932 3943
rect 2420 3937 2524 3943
rect 2692 3937 2732 3943
rect 2740 3937 3164 3943
rect 3172 3937 4348 3943
rect 4404 3937 4652 3943
rect 4660 3937 4956 3943
rect 4996 3937 5164 3943
rect 5172 3937 5260 3943
rect 5348 3937 5372 3943
rect 5492 3937 5852 3943
rect 5876 3937 5948 3943
rect 6868 3937 6908 3943
rect 6916 3937 7292 3943
rect 7300 3937 7452 3943
rect 7684 3937 7932 3943
rect 644 3917 780 3923
rect 788 3917 844 3923
rect 1220 3917 1388 3923
rect 1588 3917 1628 3923
rect 1876 3917 1884 3923
rect 2436 3917 2508 3923
rect 2564 3917 2668 3923
rect 2708 3917 2732 3923
rect 2964 3917 3148 3923
rect 3316 3917 3612 3923
rect 3636 3917 3692 3923
rect 3716 3917 3740 3923
rect 3764 3917 3788 3923
rect 3828 3917 5452 3923
rect 5524 3917 5708 3923
rect 5748 3917 5804 3923
rect 5844 3917 6236 3923
rect 6564 3917 6876 3923
rect 6916 3917 7084 3923
rect 7684 3917 7708 3923
rect 7956 3917 8060 3923
rect 36 3897 92 3903
rect 212 3897 236 3903
rect 420 3897 556 3903
rect 676 3897 780 3903
rect 788 3897 812 3903
rect 820 3897 844 3903
rect 852 3897 876 3903
rect 1524 3897 1628 3903
rect 1764 3897 1804 3903
rect 1908 3897 1964 3903
rect 2100 3897 2284 3903
rect 2356 3897 3180 3903
rect 3188 3897 3452 3903
rect 3460 3897 3484 3903
rect 3492 3897 3516 3903
rect 3540 3897 3708 3903
rect 3732 3897 3763 3903
rect 724 3877 892 3883
rect 900 3877 1004 3883
rect 1012 3877 1052 3883
rect 1108 3877 1148 3883
rect 1316 3877 1452 3883
rect 1460 3877 1964 3883
rect 1972 3877 2044 3883
rect 2308 3877 2460 3883
rect 2644 3877 2684 3883
rect 2740 3877 2780 3883
rect 2836 3877 2956 3883
rect 2980 3877 3052 3883
rect 3220 3877 3436 3883
rect 3492 3877 3548 3883
rect 3588 3877 3628 3883
rect 3716 3877 3724 3883
rect 3757 3883 3763 3897
rect 3780 3897 3852 3903
rect 3892 3897 4060 3903
rect 4084 3897 4204 3903
rect 4340 3897 5180 3903
rect 5204 3897 5228 3903
rect 5268 3897 5404 3903
rect 5412 3897 5644 3903
rect 5700 3897 5740 3903
rect 5764 3897 5932 3903
rect 5940 3897 5948 3903
rect 5956 3897 5996 3903
rect 6036 3897 6060 3903
rect 6228 3897 6396 3903
rect 6500 3897 6588 3903
rect 6676 3897 6732 3903
rect 6868 3897 6908 3903
rect 7332 3897 7356 3903
rect 7380 3897 7468 3903
rect 7572 3897 7708 3903
rect 7876 3897 7948 3903
rect 7972 3897 8044 3903
rect 8052 3897 8092 3903
rect 3757 3877 3980 3883
rect 4116 3877 4476 3883
rect 4580 3877 5132 3883
rect 5140 3877 5292 3883
rect 5316 3877 5452 3883
rect 5645 3883 5651 3896
rect 5645 3877 5788 3883
rect 5796 3877 5900 3883
rect 5908 3877 5980 3883
rect 5988 3877 6236 3883
rect 6628 3877 6716 3883
rect 6804 3877 6892 3883
rect 6900 3877 7132 3883
rect 7140 3877 7164 3883
rect 7300 3877 7388 3883
rect 7540 3877 7980 3883
rect 532 3857 684 3863
rect 868 3857 1020 3863
rect 1204 3857 1356 3863
rect 1668 3857 1852 3863
rect 1892 3857 1916 3863
rect 2020 3857 2092 3863
rect 2452 3857 2572 3863
rect 2612 3857 2700 3863
rect 2740 3857 2796 3863
rect 2836 3857 2924 3863
rect 3012 3857 3052 3863
rect 3060 3857 3116 3863
rect 3156 3857 3315 3863
rect 36 3837 220 3843
rect 500 3837 1244 3843
rect 1268 3837 1836 3843
rect 2804 3837 2908 3843
rect 2932 3837 3244 3843
rect 3252 3837 3276 3843
rect 3309 3843 3315 3857
rect 3348 3857 3452 3863
rect 3460 3857 3564 3863
rect 3572 3857 3596 3863
rect 3620 3857 3740 3863
rect 3796 3857 4028 3863
rect 4036 3857 4172 3863
rect 4804 3857 4876 3863
rect 5300 3857 5420 3863
rect 5636 3857 5756 3863
rect 5860 3857 5900 3863
rect 6068 3857 6364 3863
rect 7204 3857 7260 3863
rect 7268 3857 7404 3863
rect 7732 3857 7756 3863
rect 7908 3857 7939 3863
rect 3309 3837 3580 3843
rect 3716 3837 3836 3843
rect 3908 3837 4140 3843
rect 4148 3837 4332 3843
rect 4548 3837 4636 3843
rect 4692 3837 4924 3843
rect 4948 3837 4956 3843
rect 4964 3837 5811 3843
rect 596 3817 668 3823
rect 676 3817 828 3823
rect 836 3817 908 3823
rect 916 3817 1036 3823
rect 1348 3817 1468 3823
rect 1476 3817 1820 3823
rect 2260 3817 3148 3823
rect 3428 3817 3532 3823
rect 3556 3817 4092 3823
rect 4212 3817 4540 3823
rect 4884 3817 4892 3823
rect 4980 3817 5052 3823
rect 5060 3817 5788 3823
rect 5805 3823 5811 3837
rect 5892 3837 6060 3843
rect 6077 3837 6908 3843
rect 6077 3823 6083 3837
rect 7933 3843 7939 3857
rect 7956 3857 8060 3863
rect 7933 3837 8012 3843
rect 5805 3817 6083 3823
rect 6580 3817 6636 3823
rect 3272 3814 3320 3816
rect 3272 3806 3276 3814
rect 3286 3806 3292 3814
rect 3300 3806 3306 3814
rect 3316 3806 3320 3814
rect 3272 3804 3320 3806
rect 6344 3814 6392 3816
rect 6344 3806 6348 3814
rect 6358 3806 6364 3814
rect 6372 3806 6378 3814
rect 6388 3806 6392 3814
rect 6344 3804 6392 3806
rect 868 3797 892 3803
rect 1300 3797 1436 3803
rect 1444 3797 1516 3803
rect 2756 3797 2844 3803
rect 2868 3797 2940 3803
rect 2948 3797 3036 3803
rect 3357 3797 4396 3803
rect 708 3777 764 3783
rect 980 3777 1068 3783
rect 3357 3783 3363 3797
rect 4404 3797 4428 3803
rect 4564 3797 4620 3803
rect 4788 3797 5763 3803
rect 2468 3777 3363 3783
rect 3380 3777 3548 3783
rect 3556 3777 3724 3783
rect 3748 3777 4412 3783
rect 4420 3777 4540 3783
rect 4708 3777 4972 3783
rect 5396 3777 5468 3783
rect 5757 3783 5763 3797
rect 5876 3797 5932 3803
rect 6084 3797 6140 3803
rect 6628 3797 6684 3803
rect 5757 3777 6428 3783
rect 8116 3777 8124 3783
rect 212 3757 1020 3763
rect 1076 3757 1276 3763
rect 1716 3757 1740 3763
rect 1748 3757 1884 3763
rect 1892 3757 2012 3763
rect 2148 3757 2220 3763
rect 2276 3757 2316 3763
rect 2404 3757 2508 3763
rect 2516 3757 2844 3763
rect 3444 3757 3468 3763
rect 3572 3757 3612 3763
rect 3636 3757 3660 3763
rect 3684 3757 3756 3763
rect 4020 3757 4204 3763
rect 4228 3757 4300 3763
rect 4580 3757 4652 3763
rect 4724 3757 4748 3763
rect 5108 3757 5260 3763
rect 5268 3757 5308 3763
rect 5332 3757 5420 3763
rect 5460 3757 5500 3763
rect 5540 3757 6012 3763
rect 6020 3757 6492 3763
rect 7044 3757 7180 3763
rect 7188 3757 7372 3763
rect 7540 3757 7660 3763
rect 7812 3757 7868 3763
rect 132 3737 316 3743
rect 548 3737 572 3743
rect 660 3737 716 3743
rect 868 3737 924 3743
rect 964 3737 988 3743
rect 1044 3737 1116 3743
rect 1492 3737 1532 3743
rect 1652 3737 1724 3743
rect 1812 3737 1900 3743
rect 2036 3737 2108 3743
rect 2116 3737 2156 3743
rect 2244 3737 2284 3743
rect 2292 3737 2604 3743
rect 2660 3737 2684 3743
rect 2692 3737 2908 3743
rect 2916 3737 2988 3743
rect 2996 3737 3196 3743
rect 3284 3737 3404 3743
rect 3412 3737 3468 3743
rect 3524 3737 3788 3743
rect 3956 3737 4076 3743
rect 4420 3737 4620 3743
rect 4996 3737 5068 3743
rect 5860 3737 5955 3743
rect 292 3717 492 3723
rect 573 3723 579 3736
rect 573 3717 700 3723
rect 724 3717 892 3723
rect 1060 3717 1084 3723
rect 1540 3717 1612 3723
rect 1828 3717 1868 3723
rect 1940 3717 1964 3723
rect 2100 3717 2140 3723
rect 2388 3717 2460 3723
rect 2484 3717 2556 3723
rect 2692 3717 2812 3723
rect 2996 3717 3052 3723
rect 3197 3723 3203 3736
rect 3197 3717 3340 3723
rect 3364 3717 3436 3723
rect 3588 3717 3628 3723
rect 3652 3717 3708 3723
rect 3716 3717 3916 3723
rect 3924 3717 4780 3723
rect 4836 3717 4924 3723
rect 5204 3717 5612 3723
rect 5796 3717 5916 3723
rect 5949 3723 5955 3737
rect 5988 3737 6156 3743
rect 6308 3737 6412 3743
rect 6436 3737 6508 3743
rect 6756 3737 6876 3743
rect 6884 3737 7020 3743
rect 7316 3737 7436 3743
rect 7460 3737 7548 3743
rect 7604 3737 7644 3743
rect 7652 3737 7836 3743
rect 7844 3737 8108 3743
rect 5949 3717 6028 3723
rect 6052 3717 6108 3723
rect 6116 3717 6156 3723
rect 6452 3717 6492 3723
rect 6628 3717 6636 3723
rect 6740 3717 6812 3723
rect 6820 3717 6860 3723
rect 6948 3717 7468 3723
rect 7476 3717 7644 3723
rect 7652 3717 7756 3723
rect 7796 3717 7820 3723
rect 7924 3717 7964 3723
rect 8052 3717 8092 3723
rect 8116 3717 8156 3723
rect 276 3697 348 3703
rect 468 3697 1116 3703
rect 1124 3697 1212 3703
rect 1588 3697 1676 3703
rect 2228 3697 2252 3703
rect 2356 3697 2396 3703
rect 2452 3697 2780 3703
rect 2788 3697 4332 3703
rect 4564 3697 4572 3703
rect 4644 3697 4668 3703
rect 4772 3697 4892 3703
rect 5796 3697 5820 3703
rect 5844 3697 6316 3703
rect 6324 3697 6588 3703
rect 6596 3697 6892 3703
rect 6900 3697 6988 3703
rect 7140 3697 7148 3703
rect 7156 3697 7340 3703
rect 7348 3697 7484 3703
rect 7508 3697 7612 3703
rect 7917 3703 7923 3716
rect 7636 3697 7923 3703
rect 500 3677 908 3683
rect 980 3677 1100 3683
rect 1108 3677 1244 3683
rect 1252 3677 1820 3683
rect 2900 3677 2956 3683
rect 3204 3677 3708 3683
rect 4612 3677 5740 3683
rect 5748 3677 5948 3683
rect 5972 3677 6124 3683
rect 6276 3677 6284 3683
rect 6292 3677 6524 3683
rect 6580 3677 6684 3683
rect 7124 3677 7164 3683
rect 7428 3677 7900 3683
rect 772 3657 812 3663
rect 1524 3657 1548 3663
rect 1556 3657 1660 3663
rect 1668 3657 1724 3663
rect 3268 3657 3500 3663
rect 3940 3657 4860 3663
rect 4916 3657 4924 3663
rect 4932 3657 5020 3663
rect 5300 3657 5603 3663
rect 484 3637 1804 3643
rect 2772 3637 2796 3643
rect 3044 3637 3276 3643
rect 3460 3637 3980 3643
rect 4276 3637 4604 3643
rect 4708 3637 4732 3643
rect 4820 3637 4988 3643
rect 5556 3637 5580 3643
rect 5597 3643 5603 3657
rect 5684 3657 5788 3663
rect 5924 3657 6252 3663
rect 6628 3657 6828 3663
rect 7588 3657 7788 3663
rect 7828 3657 7852 3663
rect 5597 3637 6620 3643
rect 804 3617 940 3623
rect 1844 3617 3580 3623
rect 5444 3617 5884 3623
rect 5972 3617 6044 3623
rect 6244 3617 6652 3623
rect 6660 3617 7212 3623
rect 1736 3614 1784 3616
rect 1736 3606 1740 3614
rect 1750 3606 1756 3614
rect 1764 3606 1770 3614
rect 1780 3606 1784 3614
rect 1736 3604 1784 3606
rect 4808 3614 4856 3616
rect 4808 3606 4812 3614
rect 4822 3606 4828 3614
rect 4836 3606 4842 3614
rect 4852 3606 4856 3614
rect 4808 3604 4856 3606
rect 420 3597 572 3603
rect 3972 3597 4300 3603
rect 4340 3597 4636 3603
rect 4644 3597 4748 3603
rect 5348 3597 5372 3603
rect 5444 3597 5500 3603
rect 5940 3597 5980 3603
rect 6036 3597 6284 3603
rect 1140 3577 1452 3583
rect 2324 3577 2396 3583
rect 2404 3577 2620 3583
rect 2628 3577 2796 3583
rect 2916 3577 3052 3583
rect 3060 3577 3196 3583
rect 3524 3577 4524 3583
rect 4628 3577 4940 3583
rect 5188 3577 6140 3583
rect 6180 3577 6524 3583
rect 1108 3557 1292 3563
rect 1380 3557 1516 3563
rect 2324 3557 2492 3563
rect 2500 3557 2604 3563
rect 2612 3557 2924 3563
rect 2948 3557 3436 3563
rect 3748 3557 3772 3563
rect 3812 3557 3852 3563
rect 3972 3557 4444 3563
rect 4452 3557 4684 3563
rect 4692 3557 5292 3563
rect 5348 3557 5427 3563
rect 1012 3537 1356 3543
rect 1364 3537 1404 3543
rect 1412 3537 1484 3543
rect 1492 3537 1500 3543
rect 1620 3537 1852 3543
rect 2596 3537 2652 3543
rect 2660 3537 2892 3543
rect 2932 3537 2972 3543
rect 2996 3537 3356 3543
rect 3421 3537 3628 3543
rect 3421 3524 3427 3537
rect 3636 3537 3724 3543
rect 3732 3537 3964 3543
rect 4388 3537 4508 3543
rect 4532 3537 4540 3543
rect 5380 3537 5404 3543
rect 5421 3543 5427 3557
rect 5709 3557 5788 3563
rect 5709 3543 5715 3557
rect 6093 3557 6252 3563
rect 6093 3544 6099 3557
rect 6260 3557 6284 3563
rect 6916 3557 6972 3563
rect 7012 3557 7180 3563
rect 8084 3557 8092 3563
rect 5421 3537 5715 3543
rect 5732 3537 5804 3543
rect 5908 3537 6092 3543
rect 6132 3537 6204 3543
rect 6212 3537 6380 3543
rect 6532 3537 6620 3543
rect 6708 3537 7324 3543
rect 20 3517 76 3523
rect 84 3517 188 3523
rect 276 3517 492 3523
rect 500 3517 508 3523
rect 1236 3517 1244 3523
rect 1268 3517 1436 3523
rect 1636 3517 1884 3523
rect 2164 3517 2268 3523
rect 2356 3517 2476 3523
rect 2493 3517 2556 3523
rect 228 3497 332 3503
rect 340 3497 460 3503
rect 676 3497 860 3503
rect 868 3497 1020 3503
rect 1060 3497 1180 3503
rect 1188 3497 1228 3503
rect 1316 3497 1372 3503
rect 1444 3497 1564 3503
rect 1652 3497 1676 3503
rect 2493 3503 2499 3517
rect 2628 3517 2723 3523
rect 2717 3504 2723 3517
rect 2868 3517 3004 3523
rect 3012 3517 3212 3523
rect 3396 3517 3420 3523
rect 3604 3517 3820 3523
rect 3892 3517 4252 3523
rect 4276 3517 4556 3523
rect 4564 3517 4620 3523
rect 4836 3517 4956 3523
rect 4964 3517 5004 3523
rect 5268 3517 5404 3523
rect 5428 3517 5500 3523
rect 5524 3517 5612 3523
rect 5652 3517 5772 3523
rect 5780 3517 5852 3523
rect 5924 3517 5996 3523
rect 6068 3517 6188 3523
rect 6308 3517 6332 3523
rect 6340 3517 6476 3523
rect 6516 3517 6604 3523
rect 7156 3517 7244 3523
rect 7572 3517 7596 3523
rect 7604 3517 7724 3523
rect 7780 3517 7900 3523
rect 2276 3497 2499 3503
rect 2548 3497 2668 3503
rect 3252 3497 3356 3503
rect 3364 3497 3516 3503
rect 3780 3497 4140 3503
rect 4164 3497 4364 3503
rect 4404 3497 4444 3503
rect 4452 3497 4588 3503
rect 4596 3497 4700 3503
rect 4804 3497 4892 3503
rect 4900 3497 5036 3503
rect 5044 3497 5148 3503
rect 5204 3497 5228 3503
rect 5300 3497 5340 3503
rect 5412 3497 5452 3503
rect 5460 3497 5484 3503
rect 5492 3497 5516 3503
rect 5556 3497 5756 3503
rect 5908 3497 6236 3503
rect 6276 3497 6364 3503
rect 6372 3497 6444 3503
rect 6500 3497 6524 3503
rect 6612 3497 6716 3503
rect 6836 3497 6876 3503
rect 6884 3497 6924 3503
rect 6964 3497 7084 3503
rect 7492 3497 7516 3503
rect 7780 3497 7804 3503
rect 7812 3497 8044 3503
rect 68 3477 140 3483
rect 148 3477 380 3483
rect 548 3477 636 3483
rect 1012 3477 1340 3483
rect 1348 3477 1548 3483
rect 1556 3477 1676 3483
rect 2308 3477 2444 3483
rect 2564 3477 2604 3483
rect 2900 3477 3020 3483
rect 3140 3477 3356 3483
rect 3636 3477 3852 3483
rect 3876 3477 3996 3483
rect 4068 3477 4108 3483
rect 4372 3477 4492 3483
rect 4548 3477 4556 3483
rect 4644 3477 4812 3483
rect 5108 3477 5276 3483
rect 5284 3477 5372 3483
rect 5380 3477 5692 3483
rect 5988 3477 6540 3483
rect 6884 3477 7164 3483
rect 7396 3477 7644 3483
rect 7652 3477 7980 3483
rect 52 3457 140 3463
rect 244 3457 316 3463
rect 372 3457 476 3463
rect 1124 3457 1164 3463
rect 1172 3457 1420 3463
rect 1428 3457 1596 3463
rect 1604 3457 1708 3463
rect 2100 3457 2220 3463
rect 2484 3457 2748 3463
rect 2756 3457 3004 3463
rect 3268 3457 3388 3463
rect 3396 3457 3660 3463
rect 3668 3457 3676 3463
rect 3684 3457 3932 3463
rect 3940 3457 4028 3463
rect 4756 3457 5036 3463
rect 5044 3457 5084 3463
rect 5220 3457 5324 3463
rect 5348 3457 5420 3463
rect 5428 3457 5484 3463
rect 5524 3457 5580 3463
rect 5588 3457 5772 3463
rect 5828 3457 6060 3463
rect 6068 3457 6076 3463
rect 6100 3457 6156 3463
rect 6244 3457 6332 3463
rect 6500 3457 6700 3463
rect 7060 3457 7436 3463
rect 7668 3457 7692 3463
rect 116 3437 236 3443
rect 516 3437 540 3443
rect 932 3437 956 3443
rect 964 3437 2012 3443
rect 2676 3437 2764 3443
rect 3348 3437 3468 3443
rect 3508 3437 3564 3443
rect 3572 3437 3676 3443
rect 3684 3437 3740 3443
rect 3764 3437 3804 3443
rect 4436 3437 4796 3443
rect 4916 3437 4956 3443
rect 4980 3437 5052 3443
rect 5476 3437 5676 3443
rect 6052 3437 6124 3443
rect 6532 3437 6572 3443
rect 6804 3437 6972 3443
rect 7556 3437 7980 3443
rect 500 3417 524 3423
rect 1252 3417 1324 3423
rect 1332 3417 1740 3423
rect 1988 3417 2012 3423
rect 2756 3417 2844 3423
rect 3444 3417 3644 3423
rect 3652 3417 3692 3423
rect 3700 3417 3868 3423
rect 4676 3417 4828 3423
rect 5204 3417 5356 3423
rect 5364 3417 5404 3423
rect 5412 3417 5500 3423
rect 5508 3417 5660 3423
rect 5860 3417 5900 3423
rect 6116 3417 6188 3423
rect 6676 3417 6812 3423
rect 6820 3417 6876 3423
rect 6884 3417 7020 3423
rect 7028 3417 7068 3423
rect 3272 3414 3320 3416
rect 3272 3406 3276 3414
rect 3286 3406 3292 3414
rect 3300 3406 3306 3414
rect 3316 3406 3320 3414
rect 3272 3404 3320 3406
rect 6344 3414 6392 3416
rect 6344 3406 6348 3414
rect 6358 3406 6364 3414
rect 6372 3406 6378 3414
rect 6388 3406 6392 3414
rect 6344 3404 6392 3406
rect 740 3397 796 3403
rect 1236 3397 1612 3403
rect 1796 3397 1948 3403
rect 2436 3397 2940 3403
rect 3364 3397 3996 3403
rect 4692 3397 4748 3403
rect 5156 3397 5260 3403
rect 5332 3397 5436 3403
rect 6429 3397 7100 3403
rect 404 3377 412 3383
rect 1156 3377 1228 3383
rect 1332 3377 1836 3383
rect 1940 3377 2172 3383
rect 2484 3377 2748 3383
rect 2804 3377 2876 3383
rect 3348 3377 3388 3383
rect 3508 3377 3564 3383
rect 3620 3377 3788 3383
rect 3812 3377 3916 3383
rect 4164 3377 4204 3383
rect 4628 3377 4956 3383
rect 4964 3377 5100 3383
rect 5108 3377 5180 3383
rect 5364 3377 5468 3383
rect 5476 3377 5580 3383
rect 5588 3377 5612 3383
rect 5716 3377 5884 3383
rect 6429 3383 6435 3397
rect 7684 3397 7708 3403
rect 7716 3397 7788 3403
rect 6068 3377 6435 3383
rect 6452 3377 6588 3383
rect 6660 3377 6780 3383
rect 6788 3377 6908 3383
rect 6980 3377 7036 3383
rect 7076 3377 7132 3383
rect 7764 3377 7772 3383
rect 244 3357 396 3363
rect 740 3357 1036 3363
rect 1492 3357 1900 3363
rect 2516 3357 2588 3363
rect 2644 3357 2700 3363
rect 2772 3357 2995 3363
rect 2989 3344 2995 3357
rect 3380 3357 3420 3363
rect 3508 3357 3708 3363
rect 3828 3357 3852 3363
rect 3860 3357 4060 3363
rect 4077 3357 4172 3363
rect 84 3337 172 3343
rect 180 3337 252 3343
rect 260 3337 444 3343
rect 468 3337 572 3343
rect 644 3337 700 3343
rect 733 3337 892 3343
rect 733 3324 739 3337
rect 1732 3337 1756 3343
rect 1876 3337 2044 3343
rect 2148 3337 2204 3343
rect 2452 3337 2492 3343
rect 2548 3337 2604 3343
rect 2612 3337 2684 3343
rect 2932 3337 2956 3343
rect 2964 3337 2972 3343
rect 2996 3337 3100 3343
rect 3108 3337 3196 3343
rect 3540 3337 3660 3343
rect 3684 3337 3900 3343
rect 3908 3337 3916 3343
rect 4077 3343 4083 3357
rect 4484 3357 4716 3363
rect 4724 3357 4940 3363
rect 4948 3357 5004 3363
rect 5028 3357 5324 3363
rect 5444 3357 5596 3363
rect 5604 3357 5708 3363
rect 6084 3357 6396 3363
rect 6708 3357 6748 3363
rect 7092 3357 7212 3363
rect 7732 3357 7836 3363
rect 7844 3357 7948 3363
rect 4020 3337 4083 3343
rect 4132 3337 4236 3343
rect 4308 3337 4348 3343
rect 4628 3337 4636 3343
rect 4820 3337 4892 3343
rect 5092 3337 5148 3343
rect 5172 3337 5228 3343
rect 5508 3337 5548 3343
rect 5908 3337 6012 3343
rect 6548 3337 6652 3343
rect 6900 3337 6908 3343
rect 7460 3337 7500 3343
rect 7524 3337 7667 3343
rect 196 3317 348 3323
rect 404 3317 428 3323
rect 548 3317 604 3323
rect 692 3317 732 3323
rect 772 3317 828 3323
rect 900 3317 988 3323
rect 1076 3317 1132 3323
rect 1316 3317 3260 3323
rect 3492 3317 3756 3323
rect 3764 3317 3916 3323
rect 3924 3317 4204 3323
rect 4372 3317 4460 3323
rect 4612 3317 4732 3323
rect 4788 3317 5084 3323
rect 5140 3317 5292 3323
rect 5412 3317 5500 3323
rect 5668 3317 5788 3323
rect 6340 3317 6764 3323
rect 6868 3317 7020 3323
rect 7508 3317 7532 3323
rect 7556 3317 7612 3323
rect 7661 3323 7667 3337
rect 7684 3337 7852 3343
rect 8164 3337 8195 3343
rect 7661 3317 7740 3323
rect 7892 3317 7996 3323
rect 148 3297 204 3303
rect 436 3297 460 3303
rect 500 3297 588 3303
rect 893 3303 899 3316
rect 596 3297 899 3303
rect 1028 3297 1100 3303
rect 1492 3297 1660 3303
rect 2260 3297 2428 3303
rect 2548 3297 2652 3303
rect 2756 3297 2796 3303
rect 2884 3297 3116 3303
rect 3172 3297 3356 3303
rect 3364 3297 3628 3303
rect 3636 3297 3916 3303
rect 3988 3297 4060 3303
rect 4196 3297 4252 3303
rect 4285 3303 4291 3316
rect 4285 3297 4972 3303
rect 4980 3297 5164 3303
rect 5220 3297 5884 3303
rect 6308 3297 6364 3303
rect 7268 3297 7516 3303
rect 7604 3297 7612 3303
rect 7620 3297 7692 3303
rect 7716 3297 7756 3303
rect 7780 3297 7964 3303
rect 8036 3297 8108 3303
rect 8173 3297 8195 3303
rect 52 3277 284 3283
rect 532 3277 780 3283
rect 964 3277 1036 3283
rect 1588 3277 1612 3283
rect 1636 3277 1676 3283
rect 2468 3277 2492 3283
rect 2676 3277 3372 3283
rect 3428 3277 3612 3283
rect 3716 3277 3836 3283
rect 4740 3277 5052 3283
rect 5092 3277 5228 3283
rect 5572 3277 5740 3283
rect 5748 3277 5820 3283
rect 6132 3277 7164 3283
rect 7428 3277 7532 3283
rect 7668 3277 7692 3283
rect 7828 3277 7852 3283
rect 8173 3283 8179 3297
rect 8100 3277 8179 3283
rect 676 3257 700 3263
rect 708 3257 748 3263
rect 756 3257 940 3263
rect 1540 3257 1884 3263
rect 1892 3257 2012 3263
rect 4212 3257 4988 3263
rect 5796 3257 5932 3263
rect 6036 3257 7292 3263
rect 7636 3257 7804 3263
rect 724 3237 748 3243
rect 756 3237 1004 3243
rect 1540 3237 1612 3243
rect 1988 3237 2012 3243
rect 2116 3237 2364 3243
rect 2372 3237 2620 3243
rect 2788 3237 2812 3243
rect 4532 3237 4780 3243
rect 5060 3237 6028 3243
rect 612 3217 764 3223
rect 772 3217 924 3223
rect 1364 3217 1596 3223
rect 1892 3217 3340 3223
rect 5956 3217 5964 3223
rect 5972 3217 6108 3223
rect 6116 3217 6236 3223
rect 6244 3217 6556 3223
rect 7732 3217 7788 3223
rect 1736 3214 1784 3216
rect 1736 3206 1740 3214
rect 1750 3206 1756 3214
rect 1764 3206 1770 3214
rect 1780 3206 1784 3214
rect 1736 3204 1784 3206
rect 4808 3214 4856 3216
rect 4808 3206 4812 3214
rect 4822 3206 4828 3214
rect 4836 3206 4842 3214
rect 4852 3206 4856 3214
rect 4808 3204 4856 3206
rect 628 3197 732 3203
rect 852 3197 1068 3203
rect 1812 3197 2908 3203
rect 2916 3197 2940 3203
rect 3780 3197 4204 3203
rect 6180 3197 6268 3203
rect 6276 3197 6508 3203
rect 7092 3197 7116 3203
rect 548 3177 636 3183
rect 4068 3177 4252 3183
rect 4500 3177 4764 3183
rect 4884 3177 4892 3183
rect 5268 3177 5324 3183
rect 6244 3177 6460 3183
rect 6756 3177 6876 3183
rect 7492 3177 7516 3183
rect 7956 3177 8012 3183
rect 532 3157 668 3163
rect 1060 3157 1084 3163
rect 1092 3157 1276 3163
rect 2420 3157 2476 3163
rect 2484 3157 2556 3163
rect 2564 3157 2684 3163
rect 2692 3157 2796 3163
rect 3540 3157 3788 3163
rect 4468 3157 4604 3163
rect 4612 3157 4716 3163
rect 6420 3157 6444 3163
rect 6452 3157 6748 3163
rect 6868 3157 6972 3163
rect 6996 3157 7036 3163
rect 7460 3157 7484 3163
rect 7492 3157 7836 3163
rect 7844 3157 8028 3163
rect 484 3137 540 3143
rect 708 3137 780 3143
rect 1284 3137 1356 3143
rect 1412 3137 1436 3143
rect 1444 3137 1747 3143
rect 1741 3124 1747 3137
rect 2308 3137 2412 3143
rect 2420 3137 2460 3143
rect 3332 3137 3452 3143
rect 3476 3137 3580 3143
rect 3620 3137 3644 3143
rect 3652 3137 3692 3143
rect 3700 3137 3884 3143
rect 4516 3137 4636 3143
rect 4644 3137 4684 3143
rect 5172 3137 5932 3143
rect 5940 3137 6124 3143
rect 6324 3137 6508 3143
rect 6724 3137 7228 3143
rect 7796 3137 7932 3143
rect 100 3117 236 3123
rect 244 3117 380 3123
rect 500 3117 572 3123
rect 772 3117 828 3123
rect 1348 3117 1372 3123
rect 1572 3117 1644 3123
rect 1748 3117 1827 3123
rect 1821 3104 1827 3117
rect 1844 3117 1996 3123
rect 2196 3117 2364 3123
rect 2452 3117 2508 3123
rect 2516 3117 2652 3123
rect 2772 3117 2828 3123
rect 3428 3117 3500 3123
rect 3508 3117 3564 3123
rect 3652 3117 3740 3123
rect 3860 3117 3980 3123
rect 4420 3117 4524 3123
rect 4532 3117 4572 3123
rect 4580 3117 4652 3123
rect 4660 3117 4732 3123
rect 5140 3117 5196 3123
rect 5204 3117 5356 3123
rect 5412 3117 5484 3123
rect 5492 3117 5852 3123
rect 6148 3117 6236 3123
rect 6468 3117 6652 3123
rect 6676 3117 6860 3123
rect 6868 3117 6908 3123
rect 6948 3117 7139 3123
rect 7133 3104 7139 3117
rect 7508 3117 7532 3123
rect 7540 3117 7612 3123
rect 7812 3117 7868 3123
rect 7908 3117 8028 3123
rect 84 3097 140 3103
rect 324 3097 1004 3103
rect 1156 3097 1180 3103
rect 1348 3097 1420 3103
rect 1540 3097 1580 3103
rect 1588 3097 1660 3103
rect 1668 3097 1756 3103
rect 1828 3097 1923 3103
rect 1917 3084 1923 3097
rect 1972 3097 1980 3103
rect 1988 3097 2012 3103
rect 2500 3097 2572 3103
rect 2660 3097 2716 3103
rect 2724 3097 2780 3103
rect 3060 3097 3164 3103
rect 3188 3097 4812 3103
rect 4820 3097 4956 3103
rect 4964 3097 4988 3103
rect 5076 3097 5116 3103
rect 5684 3097 5708 3103
rect 5716 3097 5756 3103
rect 5924 3097 6012 3103
rect 6084 3097 6172 3103
rect 6324 3097 6396 3103
rect 6436 3097 6588 3103
rect 6596 3097 6716 3103
rect 6788 3097 6844 3103
rect 6980 3097 7052 3103
rect 7140 3097 7180 3103
rect 7268 3097 7292 3103
rect 7588 3097 7628 3103
rect 7636 3097 7660 3103
rect 7748 3097 7772 3103
rect 7876 3097 8012 3103
rect 8068 3097 8140 3103
rect 68 3077 108 3083
rect 164 3077 284 3083
rect 420 3077 524 3083
rect 660 3077 732 3083
rect 836 3077 892 3083
rect 916 3077 956 3083
rect 1156 3077 1203 3083
rect 20 3057 60 3063
rect 68 3057 172 3063
rect 564 3057 636 3063
rect 724 3057 764 3063
rect 1197 3063 1203 3077
rect 1220 3077 1276 3083
rect 1380 3077 1516 3083
rect 1524 3077 1724 3083
rect 1732 3077 1884 3083
rect 1924 3077 1980 3083
rect 2036 3077 2172 3083
rect 2180 3077 2316 3083
rect 2324 3077 2412 3083
rect 2468 3077 2572 3083
rect 2580 3077 2620 3083
rect 2932 3077 3132 3083
rect 3204 3077 3420 3083
rect 3460 3077 3628 3083
rect 3796 3077 3836 3083
rect 4052 3077 4076 3083
rect 4084 3077 4236 3083
rect 4420 3077 4444 3083
rect 4548 3077 4700 3083
rect 4708 3077 4956 3083
rect 5124 3077 5196 3083
rect 5348 3077 5660 3083
rect 5668 3077 5900 3083
rect 6164 3077 6220 3083
rect 6637 3077 7004 3083
rect 6637 3064 6643 3077
rect 7012 3077 7180 3083
rect 7188 3077 7228 3083
rect 7300 3077 7596 3083
rect 7604 3077 7644 3083
rect 7876 3077 8060 3083
rect 1197 3057 1388 3063
rect 1396 3057 1500 3063
rect 1508 3057 1612 3063
rect 1620 3057 1932 3063
rect 2596 3057 2652 3063
rect 3028 3057 3036 3063
rect 3348 3057 3516 3063
rect 3524 3057 3548 3063
rect 3732 3057 3804 3063
rect 3860 3057 3884 3063
rect 4340 3057 4412 3063
rect 4436 3057 4524 3063
rect 4532 3057 4556 3063
rect 4564 3057 4636 3063
rect 4676 3057 4924 3063
rect 4932 3057 4972 3063
rect 5572 3057 5724 3063
rect 6404 3057 6636 3063
rect 6660 3057 6796 3063
rect 6948 3057 6988 3063
rect 7060 3057 7340 3063
rect 7460 3057 7548 3063
rect 7572 3057 7916 3063
rect 68 3037 92 3043
rect 100 3037 188 3043
rect 436 3037 684 3043
rect 692 3037 844 3043
rect 1172 3037 1356 3043
rect 2612 3037 2652 3043
rect 2660 3037 2892 3043
rect 2900 3037 4060 3043
rect 4644 3037 4668 3043
rect 4948 3037 5068 3043
rect 5540 3037 5564 3043
rect 5572 3037 5836 3043
rect 5956 3037 6012 3043
rect 6020 3037 6140 3043
rect 6989 3043 6995 3056
rect 6724 3037 7148 3043
rect 7636 3037 7788 3043
rect 3556 3017 3772 3023
rect 3780 3017 3884 3023
rect 4404 3017 4540 3023
rect 4916 3017 4972 3023
rect 6692 3017 6764 3023
rect 6884 3017 6988 3023
rect 6996 3017 7036 3023
rect 7044 3017 7132 3023
rect 7716 3017 7772 3023
rect 3272 3014 3320 3016
rect 3272 3006 3276 3014
rect 3286 3006 3292 3014
rect 3300 3006 3306 3014
rect 3316 3006 3320 3014
rect 3272 3004 3320 3006
rect 6344 3014 6392 3016
rect 6344 3006 6348 3014
rect 6358 3006 6364 3014
rect 6372 3006 6378 3014
rect 6388 3006 6392 3014
rect 6344 3004 6392 3006
rect 468 2997 556 3003
rect 1012 2997 1324 3003
rect 1412 2997 1564 3003
rect 1572 2997 1708 3003
rect 3476 2997 3532 3003
rect 3908 2997 4044 3003
rect 5492 2997 5596 3003
rect 5668 2997 5804 3003
rect 5844 2997 5996 3003
rect 6436 2997 6732 3003
rect 6852 2997 6924 3003
rect 6980 2997 7420 3003
rect 7428 2997 7516 3003
rect 7524 2997 7676 3003
rect 7684 2997 7724 3003
rect 564 2977 620 2983
rect 628 2977 796 2983
rect 1268 2977 1324 2983
rect 1332 2977 1724 2983
rect 1732 2977 1836 2983
rect 2020 2977 2332 2983
rect 2340 2977 2380 2983
rect 2468 2977 2492 2983
rect 2500 2977 2572 2983
rect 2996 2977 3180 2983
rect 3380 2977 3484 2983
rect 3508 2977 3532 2983
rect 3540 2977 3644 2983
rect 3652 2977 3676 2983
rect 3684 2977 3756 2983
rect 3764 2977 4172 2983
rect 5268 2977 5388 2983
rect 5396 2977 5468 2983
rect 5572 2977 6348 2983
rect 6356 2977 6540 2983
rect 6852 2977 6956 2983
rect 7716 2977 7836 2983
rect 372 2957 828 2963
rect 836 2957 988 2963
rect 996 2957 1132 2963
rect 1700 2957 2044 2963
rect 2100 2957 2220 2963
rect 2500 2957 2620 2963
rect 3156 2957 3356 2963
rect 3412 2957 3644 2963
rect 3652 2957 3660 2963
rect 3668 2957 3772 2963
rect 3780 2957 3980 2963
rect 4292 2957 4460 2963
rect 4548 2957 4588 2963
rect 5540 2957 5612 2963
rect 6580 2957 6636 2963
rect 6644 2957 6892 2963
rect 6916 2957 7372 2963
rect 7380 2957 7388 2963
rect 7444 2957 7500 2963
rect 7668 2957 7932 2963
rect 36 2937 60 2943
rect 148 2937 188 2943
rect 228 2937 300 2943
rect 500 2937 588 2943
rect 788 2937 924 2943
rect 1092 2937 1164 2943
rect 1364 2937 1580 2943
rect 1588 2937 1644 2943
rect 1716 2937 1932 2943
rect 1940 2937 2028 2943
rect 2308 2937 2348 2943
rect 2356 2937 2396 2943
rect 2452 2937 2556 2943
rect 2596 2937 2940 2943
rect 3332 2937 3484 2943
rect 3524 2937 3804 2943
rect 3812 2937 3996 2943
rect 4100 2937 4236 2943
rect 4324 2937 4412 2943
rect 4436 2937 4556 2943
rect 4740 2937 4860 2943
rect 5092 2937 5148 2943
rect 5364 2937 5548 2943
rect 5716 2937 5756 2943
rect 5796 2937 5900 2943
rect 6580 2937 6620 2943
rect 6948 2937 7036 2943
rect 7364 2937 7596 2943
rect 52 2917 204 2923
rect 1444 2917 1628 2923
rect 1668 2917 1740 2923
rect 1764 2917 1948 2923
rect 2036 2917 2156 2923
rect 2468 2917 2508 2923
rect 2580 2917 2684 2923
rect 2932 2917 3052 2923
rect 3204 2917 3388 2923
rect 3460 2917 3628 2923
rect 3636 2917 3644 2923
rect 3828 2917 3852 2923
rect 3876 2917 4140 2923
rect 4452 2917 4460 2923
rect 4468 2917 4620 2923
rect 5156 2917 5164 2923
rect 5444 2917 5580 2923
rect 5588 2917 5740 2923
rect 5828 2917 6092 2923
rect 6484 2917 6588 2923
rect 6612 2917 6700 2923
rect 6772 2917 6860 2923
rect 6932 2917 7036 2923
rect 7044 2917 7068 2923
rect 7092 2917 7132 2923
rect 7412 2917 7484 2923
rect 7748 2917 7788 2923
rect 8004 2917 8028 2923
rect 36 2897 140 2903
rect 180 2897 204 2903
rect 1860 2897 2012 2903
rect 2388 2897 2700 2903
rect 2708 2897 2892 2903
rect 2900 2897 3571 2903
rect 756 2877 812 2883
rect 820 2877 876 2883
rect 1556 2877 1612 2883
rect 1620 2877 1804 2883
rect 2532 2877 2908 2883
rect 3332 2877 3548 2883
rect 3565 2883 3571 2897
rect 3604 2897 3820 2903
rect 3828 2897 3916 2903
rect 3956 2897 3996 2903
rect 4404 2897 4444 2903
rect 4452 2897 4476 2903
rect 4516 2897 4604 2903
rect 4612 2897 4700 2903
rect 4708 2897 4796 2903
rect 4900 2897 4908 2903
rect 5076 2897 6252 2903
rect 6948 2897 7292 2903
rect 7476 2897 7628 2903
rect 7844 2897 7932 2903
rect 8164 2897 8195 2903
rect 3565 2877 5212 2883
rect 5444 2877 5660 2883
rect 6340 2877 6508 2883
rect 6516 2877 6668 2883
rect 7892 2877 7996 2883
rect 52 2857 76 2863
rect 84 2857 188 2863
rect 196 2857 364 2863
rect 372 2857 748 2863
rect 1252 2857 2108 2863
rect 2916 2857 3164 2863
rect 3428 2857 3580 2863
rect 3588 2857 4076 2863
rect 4084 2857 4124 2863
rect 4372 2857 4956 2863
rect 4964 2857 5196 2863
rect 5204 2857 5308 2863
rect 7908 2857 7932 2863
rect 740 2837 780 2843
rect 1540 2837 1548 2843
rect 2820 2837 2876 2843
rect 2884 2837 3196 2843
rect 3524 2837 3676 2843
rect 3940 2837 4124 2843
rect 4580 2837 4684 2843
rect 5060 2837 5436 2843
rect 5460 2837 5676 2843
rect 5684 2837 5756 2843
rect 4308 2817 4748 2823
rect 5284 2817 5516 2823
rect 5588 2817 5724 2823
rect 6148 2817 7148 2823
rect 1736 2814 1784 2816
rect 1736 2806 1740 2814
rect 1750 2806 1756 2814
rect 1764 2806 1770 2814
rect 1780 2806 1784 2814
rect 1736 2804 1784 2806
rect 4808 2814 4856 2816
rect 4808 2806 4812 2814
rect 4822 2806 4828 2814
rect 4836 2806 4842 2814
rect 4852 2806 4856 2814
rect 4808 2804 4856 2806
rect 2468 2797 2860 2803
rect 2868 2797 3132 2803
rect 4372 2797 4540 2803
rect 4644 2797 4700 2803
rect 5252 2797 5292 2803
rect 5300 2797 5500 2803
rect 5508 2797 5596 2803
rect 5604 2797 5708 2803
rect 5892 2797 7068 2803
rect 7076 2797 7180 2803
rect 7188 2797 7324 2803
rect 212 2777 236 2783
rect 1860 2777 2140 2783
rect 2148 2777 2300 2783
rect 2932 2777 2956 2783
rect 2964 2777 3116 2783
rect 4212 2777 4771 2783
rect 4765 2764 4771 2777
rect 4804 2777 6300 2783
rect 6308 2777 6956 2783
rect 6964 2777 6988 2783
rect 7396 2777 7484 2783
rect 7812 2777 8028 2783
rect 420 2757 508 2763
rect 1460 2757 1884 2763
rect 4244 2757 4668 2763
rect 4772 2757 5068 2763
rect 5524 2757 5692 2763
rect 7428 2757 8012 2763
rect 276 2737 396 2743
rect 964 2737 1436 2743
rect 1444 2737 1884 2743
rect 2084 2737 2108 2743
rect 3252 2737 3548 2743
rect 3556 2737 3788 2743
rect 3892 2737 4060 2743
rect 4068 2737 4508 2743
rect 4628 2737 4684 2743
rect 5364 2737 5516 2743
rect 5700 2737 5740 2743
rect 5940 2737 6108 2743
rect 6116 2737 6172 2743
rect 6276 2737 6300 2743
rect 7364 2737 7868 2743
rect 7908 2737 7964 2743
rect 164 2717 316 2723
rect 436 2717 604 2723
rect 957 2723 963 2736
rect 628 2717 963 2723
rect 1060 2717 1164 2723
rect 1428 2717 1580 2723
rect 1620 2717 1644 2723
rect 2052 2717 2364 2723
rect 3204 2717 3724 2723
rect 4276 2717 4412 2723
rect 4676 2717 4716 2723
rect 4724 2717 4780 2723
rect 4788 2717 4892 2723
rect 4900 2717 5004 2723
rect 5012 2717 5084 2723
rect 5172 2717 5324 2723
rect 5396 2717 5484 2723
rect 5524 2717 5580 2723
rect 5892 2717 5948 2723
rect 7156 2717 7404 2723
rect 7524 2717 7564 2723
rect 7940 2717 8060 2723
rect 132 2697 268 2703
rect 276 2697 492 2703
rect 500 2697 572 2703
rect 836 2697 892 2703
rect 1076 2697 1116 2703
rect 1316 2697 1628 2703
rect 1645 2697 1820 2703
rect 116 2677 428 2683
rect 612 2677 860 2683
rect 868 2677 876 2683
rect 948 2677 988 2683
rect 996 2677 1100 2683
rect 1108 2677 1132 2683
rect 1645 2683 1651 2697
rect 1844 2697 1948 2703
rect 2068 2697 2172 2703
rect 2484 2697 2524 2703
rect 2532 2697 2684 2703
rect 2804 2697 2988 2703
rect 3060 2697 3180 2703
rect 3396 2697 3452 2703
rect 3492 2697 3580 2703
rect 4500 2697 4556 2703
rect 4621 2697 4748 2703
rect 1572 2677 1651 2683
rect 1684 2677 2012 2683
rect 2132 2677 2140 2683
rect 2148 2677 2236 2683
rect 2420 2677 2620 2683
rect 2628 2677 2700 2683
rect 3108 2677 3692 2683
rect 3700 2677 3836 2683
rect 4180 2677 4220 2683
rect 4292 2677 4460 2683
rect 4621 2683 4627 2697
rect 5012 2697 5148 2703
rect 5188 2697 5260 2703
rect 5476 2697 5708 2703
rect 5860 2697 5900 2703
rect 6100 2697 6268 2703
rect 6308 2697 6636 2703
rect 6788 2697 7052 2703
rect 7220 2697 7260 2703
rect 7268 2697 7452 2703
rect 7604 2697 7804 2703
rect 7924 2697 7948 2703
rect 4564 2677 4627 2683
rect 4644 2677 4668 2683
rect 4676 2677 4732 2683
rect 5140 2677 5212 2683
rect 5412 2677 5532 2683
rect 5540 2677 5564 2683
rect 5572 2677 5756 2683
rect 5780 2677 5820 2683
rect 5892 2677 5948 2683
rect 5972 2677 5996 2683
rect 6004 2677 6508 2683
rect 6660 2677 6684 2683
rect 6692 2677 6716 2683
rect 7348 2677 7420 2683
rect 7428 2677 7484 2683
rect 7588 2677 7676 2683
rect 7860 2677 7948 2683
rect 8068 2677 8092 2683
rect 772 2657 796 2663
rect 852 2657 1020 2663
rect 1700 2657 1788 2663
rect 1956 2657 1980 2663
rect 2004 2657 2060 2663
rect 2388 2657 2732 2663
rect 3172 2657 3196 2663
rect 3252 2657 3388 2663
rect 3396 2657 3420 2663
rect 3428 2657 3596 2663
rect 3604 2657 3692 2663
rect 3764 2657 3836 2663
rect 4548 2657 4556 2663
rect 4596 2657 4652 2663
rect 5268 2657 5436 2663
rect 5556 2657 5724 2663
rect 5748 2657 5868 2663
rect 5988 2657 6012 2663
rect 6148 2657 6268 2663
rect 7380 2657 7452 2663
rect 7460 2657 7532 2663
rect 7588 2657 7836 2663
rect 7844 2657 7868 2663
rect 7876 2657 7964 2663
rect 484 2637 732 2643
rect 932 2637 2316 2643
rect 2452 2637 2492 2643
rect 2564 2637 2636 2643
rect 2964 2637 3452 2643
rect 4461 2637 4556 2643
rect 1620 2617 1820 2623
rect 1828 2617 1868 2623
rect 1876 2617 2076 2623
rect 2445 2623 2451 2636
rect 2132 2617 2451 2623
rect 2532 2617 2668 2623
rect 3460 2617 3724 2623
rect 4020 2617 4268 2623
rect 4461 2623 4467 2637
rect 4628 2637 5148 2643
rect 5188 2637 5692 2643
rect 5732 2637 5804 2643
rect 5812 2637 6140 2643
rect 6148 2637 6284 2643
rect 6292 2637 6428 2643
rect 6964 2637 7308 2643
rect 7316 2637 7388 2643
rect 7684 2637 7852 2643
rect 4324 2617 4467 2623
rect 4484 2617 4652 2623
rect 5172 2617 5612 2623
rect 5716 2617 5916 2623
rect 6756 2617 6940 2623
rect 6948 2617 7788 2623
rect 3272 2614 3320 2616
rect 3272 2606 3276 2614
rect 3286 2606 3292 2614
rect 3300 2606 3306 2614
rect 3316 2606 3320 2614
rect 3272 2604 3320 2606
rect 6344 2614 6392 2616
rect 6344 2606 6348 2614
rect 6358 2606 6364 2614
rect 6372 2606 6378 2614
rect 6388 2606 6392 2614
rect 6344 2604 6392 2606
rect 484 2597 1036 2603
rect 1508 2597 1612 2603
rect 1780 2597 2252 2603
rect 2868 2597 2972 2603
rect 2980 2597 3100 2603
rect 4100 2597 4108 2603
rect 4116 2597 4220 2603
rect 4260 2597 4604 2603
rect 4788 2597 4828 2603
rect 5572 2597 6060 2603
rect 6068 2597 6236 2603
rect 6772 2597 7516 2603
rect 7524 2597 7564 2603
rect 7572 2597 7644 2603
rect 8068 2597 8108 2603
rect 548 2577 588 2583
rect 948 2577 1292 2583
rect 1316 2577 1388 2583
rect 1396 2577 1516 2583
rect 1604 2577 1628 2583
rect 1636 2577 1660 2583
rect 1668 2577 1964 2583
rect 1988 2577 2028 2583
rect 2148 2577 2908 2583
rect 3092 2577 3244 2583
rect 3540 2577 3708 2583
rect 3716 2577 3788 2583
rect 4036 2577 4076 2583
rect 4148 2577 4204 2583
rect 4308 2577 4460 2583
rect 4468 2577 4540 2583
rect 4548 2577 4604 2583
rect 5124 2577 5308 2583
rect 5668 2577 6124 2583
rect 6132 2577 6204 2583
rect 6212 2577 6412 2583
rect 7284 2577 7468 2583
rect 8084 2577 8108 2583
rect 516 2557 540 2563
rect 804 2557 908 2563
rect 932 2557 988 2563
rect 1348 2557 1484 2563
rect 1492 2557 1772 2563
rect 1796 2557 1932 2563
rect 2068 2557 2588 2563
rect 2596 2557 2876 2563
rect 3124 2557 3228 2563
rect 3236 2557 3260 2563
rect 3268 2557 3436 2563
rect 3972 2557 4156 2563
rect 4228 2557 4444 2563
rect 4452 2557 4540 2563
rect 4580 2557 4636 2563
rect 4756 2557 4956 2563
rect 5012 2557 5324 2563
rect 5588 2557 5740 2563
rect 5764 2557 5868 2563
rect 6020 2557 6156 2563
rect 6164 2557 6252 2563
rect 6356 2557 6444 2563
rect 7124 2557 7356 2563
rect 7364 2557 7660 2563
rect 7748 2557 7916 2563
rect 148 2537 620 2543
rect 900 2537 1004 2543
rect 1012 2537 1084 2543
rect 1092 2537 1228 2543
rect 1636 2537 1692 2543
rect 1725 2537 1836 2543
rect 1725 2524 1731 2537
rect 1892 2537 2076 2543
rect 2084 2537 2124 2543
rect 2228 2537 2284 2543
rect 2292 2537 2364 2543
rect 2484 2537 2572 2543
rect 3220 2537 3308 2543
rect 3364 2537 3500 2543
rect 3604 2537 3804 2543
rect 3828 2537 3868 2543
rect 3892 2537 3932 2543
rect 3940 2537 4604 2543
rect 4692 2537 4748 2543
rect 5188 2537 5260 2543
rect 5364 2537 5484 2543
rect 5652 2537 5724 2543
rect 5860 2537 5964 2543
rect 5972 2537 6028 2543
rect 6244 2537 6524 2543
rect 6596 2537 6780 2543
rect 7085 2537 7228 2543
rect 7085 2524 7091 2537
rect 7556 2537 7884 2543
rect 820 2517 844 2523
rect 868 2517 892 2523
rect 980 2517 1036 2523
rect 1268 2517 1356 2523
rect 1364 2517 1548 2523
rect 1556 2517 1724 2523
rect 1748 2517 1852 2523
rect 1924 2517 1980 2523
rect 2260 2517 2348 2523
rect 2372 2517 2492 2523
rect 2500 2517 2540 2523
rect 2916 2517 3036 2523
rect 3044 2517 3132 2523
rect 3172 2517 3468 2523
rect 3716 2517 3900 2523
rect 4196 2517 4380 2523
rect 4404 2517 4476 2523
rect 4548 2517 5020 2523
rect 5220 2517 5404 2523
rect 5508 2517 5612 2523
rect 5620 2517 5660 2523
rect 5700 2517 5740 2523
rect 5860 2517 6108 2523
rect 6116 2517 6172 2523
rect 6260 2517 6268 2523
rect 6276 2517 6364 2523
rect 6436 2517 6620 2523
rect 6692 2517 6812 2523
rect 7220 2517 7340 2523
rect 7508 2517 7580 2523
rect 7636 2517 7676 2523
rect 7716 2517 7740 2523
rect 7812 2517 7836 2523
rect 516 2497 940 2503
rect 1028 2497 1100 2503
rect 1108 2497 1132 2503
rect 1236 2497 1260 2503
rect 1348 2497 1468 2503
rect 1524 2497 1612 2503
rect 1620 2497 2108 2503
rect 2436 2497 2684 2503
rect 2900 2497 2988 2503
rect 2996 2497 3180 2503
rect 3188 2497 3420 2503
rect 3428 2497 3484 2503
rect 3652 2497 4108 2503
rect 4116 2497 4556 2503
rect 4564 2497 5564 2503
rect 5741 2503 5747 2516
rect 5741 2497 5932 2503
rect 5940 2497 5980 2503
rect 6036 2497 6076 2503
rect 6212 2497 6268 2503
rect 7188 2497 7244 2503
rect 7748 2497 7804 2503
rect 8029 2497 8195 2503
rect 900 2477 1068 2483
rect 1076 2477 1148 2483
rect 1492 2477 1516 2483
rect 1540 2477 1692 2483
rect 1700 2477 1788 2483
rect 1844 2477 1900 2483
rect 2964 2477 3196 2483
rect 3284 2477 3356 2483
rect 3476 2477 3532 2483
rect 3588 2477 3660 2483
rect 4276 2477 4396 2483
rect 4484 2477 4620 2483
rect 4708 2477 4764 2483
rect 5380 2477 6291 2483
rect 740 2457 1276 2463
rect 1668 2457 1884 2463
rect 2804 2457 3052 2463
rect 4116 2457 4284 2463
rect 4356 2457 4428 2463
rect 4436 2457 4764 2463
rect 4772 2457 5052 2463
rect 5892 2457 5916 2463
rect 5924 2457 6220 2463
rect 6285 2463 6291 2477
rect 6308 2477 6540 2483
rect 6612 2477 6668 2483
rect 8029 2483 8035 2497
rect 7796 2477 8035 2483
rect 6285 2457 7276 2463
rect 852 2437 956 2443
rect 964 2437 1036 2443
rect 4372 2437 4428 2443
rect 4996 2437 7356 2443
rect 7364 2437 7484 2443
rect 7492 2437 7580 2443
rect 7588 2437 7612 2443
rect 4420 2417 4588 2423
rect 1736 2414 1784 2416
rect 1736 2406 1740 2414
rect 1750 2406 1756 2414
rect 1764 2406 1770 2414
rect 1780 2406 1784 2414
rect 1736 2404 1784 2406
rect 4808 2414 4856 2416
rect 4808 2406 4812 2414
rect 4822 2406 4828 2414
rect 4836 2406 4842 2414
rect 4852 2406 4856 2414
rect 4808 2404 4856 2406
rect 484 2397 572 2403
rect 1188 2397 1484 2403
rect 2324 2397 3180 2403
rect 4596 2397 4716 2403
rect 5060 2397 5132 2403
rect 5140 2397 5212 2403
rect 788 2377 844 2383
rect 852 2377 1164 2383
rect 1172 2377 1340 2383
rect 1428 2377 2060 2383
rect 2468 2377 2876 2383
rect 3172 2377 3356 2383
rect 4068 2377 4076 2383
rect 4148 2377 4300 2383
rect 4516 2377 4812 2383
rect 4820 2377 5004 2383
rect 5460 2377 5756 2383
rect 6868 2377 6972 2383
rect 7428 2377 7516 2383
rect 308 2357 364 2363
rect 516 2357 604 2363
rect 1124 2357 1548 2363
rect 1572 2357 2028 2363
rect 2644 2357 2924 2363
rect 3924 2357 3996 2363
rect 4260 2357 4764 2363
rect 4772 2357 4876 2363
rect 5396 2357 5516 2363
rect 5524 2357 5740 2363
rect 5924 2357 5980 2363
rect 6116 2357 6284 2363
rect 6676 2357 6764 2363
rect 6772 2357 6844 2363
rect 6852 2357 6924 2363
rect 7012 2357 7036 2363
rect 7348 2357 7740 2363
rect 7748 2357 7772 2363
rect 356 2337 1260 2343
rect 1268 2337 1468 2343
rect 2852 2337 2892 2343
rect 3028 2337 3276 2343
rect 4244 2337 4332 2343
rect 4404 2337 4556 2343
rect 4564 2337 4668 2343
rect 4701 2337 4940 2343
rect 4701 2324 4707 2337
rect 5652 2337 5804 2343
rect 5812 2337 5820 2343
rect 5924 2337 6124 2343
rect 6148 2337 6188 2343
rect 6468 2337 6908 2343
rect 7044 2337 7100 2343
rect 7108 2337 7228 2343
rect 7524 2337 7740 2343
rect 7812 2337 7884 2343
rect 212 2317 380 2323
rect 388 2317 444 2323
rect 452 2317 508 2323
rect 548 2317 652 2323
rect 980 2317 1052 2323
rect 1124 2317 1180 2323
rect 1188 2317 1228 2323
rect 1396 2317 1532 2323
rect 1908 2317 2236 2323
rect 2740 2317 2796 2323
rect 2804 2317 2988 2323
rect 3076 2317 3148 2323
rect 3156 2317 3964 2323
rect 4276 2317 4492 2323
rect 4532 2317 4572 2323
rect 4644 2317 4700 2323
rect 4772 2317 4780 2323
rect 4836 2317 5020 2323
rect 5028 2317 5068 2323
rect 5508 2317 5628 2323
rect 6068 2317 6204 2323
rect 6324 2317 6428 2323
rect 6804 2317 6876 2323
rect 6996 2317 7116 2323
rect 7412 2317 7564 2323
rect 7588 2317 7756 2323
rect 7764 2317 7788 2323
rect 612 2297 764 2303
rect 1060 2297 1100 2303
rect 1140 2297 1308 2303
rect 1380 2297 1436 2303
rect 1556 2297 1692 2303
rect 1876 2297 1900 2303
rect 1956 2297 2012 2303
rect 2020 2297 2060 2303
rect 2068 2297 2252 2303
rect 2628 2297 2668 2303
rect 2676 2297 2780 2303
rect 2804 2297 2844 2303
rect 2852 2297 3004 2303
rect 3348 2297 3404 2303
rect 3476 2297 3548 2303
rect 3556 2297 3708 2303
rect 3716 2297 3756 2303
rect 3812 2297 3996 2303
rect 4068 2297 4092 2303
rect 4100 2297 4252 2303
rect 4372 2297 4412 2303
rect 4452 2297 4748 2303
rect 4756 2297 4828 2303
rect 4996 2297 5084 2303
rect 5108 2297 5244 2303
rect 5412 2297 5596 2303
rect 5684 2297 5820 2303
rect 5844 2297 5923 2303
rect 116 2277 348 2283
rect 356 2277 412 2283
rect 420 2277 476 2283
rect 1140 2277 1212 2283
rect 1220 2277 1356 2283
rect 1444 2277 1596 2283
rect 1972 2277 2108 2283
rect 2116 2277 2428 2283
rect 2436 2277 2476 2283
rect 2868 2277 3036 2283
rect 3108 2277 3148 2283
rect 3732 2277 3964 2283
rect 4196 2277 5260 2283
rect 5460 2277 5516 2283
rect 5540 2277 5580 2283
rect 5636 2277 5692 2283
rect 5796 2277 5852 2283
rect 5860 2277 5900 2283
rect 5917 2283 5923 2297
rect 5940 2297 6300 2303
rect 6756 2297 6892 2303
rect 6948 2297 6988 2303
rect 6996 2297 7244 2303
rect 7252 2297 7500 2303
rect 7604 2297 7660 2303
rect 7732 2297 7788 2303
rect 7828 2297 7852 2303
rect 7924 2297 7980 2303
rect 5917 2277 6076 2283
rect 6116 2277 6172 2283
rect 6212 2277 6460 2283
rect 6468 2277 6860 2283
rect 7476 2277 7676 2283
rect 7684 2277 7852 2283
rect 7860 2277 7916 2283
rect 7924 2277 8108 2283
rect 1012 2257 1644 2263
rect 1876 2257 2092 2263
rect 2388 2257 2556 2263
rect 2580 2257 2636 2263
rect 2644 2257 2700 2263
rect 2724 2257 2835 2263
rect 196 2237 220 2243
rect 276 2237 300 2243
rect 1348 2237 1404 2243
rect 1908 2237 2092 2243
rect 2356 2237 2588 2243
rect 2644 2237 2812 2243
rect 2829 2243 2835 2257
rect 2964 2257 3052 2263
rect 3172 2257 3388 2263
rect 3828 2257 4508 2263
rect 4548 2257 4652 2263
rect 4692 2257 4780 2263
rect 4932 2257 5020 2263
rect 5604 2257 5644 2263
rect 5668 2257 5724 2263
rect 5748 2257 5916 2263
rect 5924 2257 5964 2263
rect 6260 2257 6332 2263
rect 7460 2257 7516 2263
rect 7620 2257 7836 2263
rect 2829 2237 3500 2243
rect 4388 2237 4460 2243
rect 4477 2237 4524 2243
rect 164 2217 188 2223
rect 1252 2217 2268 2223
rect 2372 2217 2572 2223
rect 2660 2217 2796 2223
rect 3540 2217 3852 2223
rect 3860 2217 4348 2223
rect 4477 2223 4483 2237
rect 4564 2237 4844 2243
rect 4900 2237 4956 2243
rect 5908 2237 6156 2243
rect 6420 2237 6540 2243
rect 6660 2237 6716 2243
rect 6740 2237 6764 2243
rect 6772 2237 6812 2243
rect 4420 2217 4483 2223
rect 4500 2217 4572 2223
rect 4660 2217 5084 2223
rect 5892 2217 6012 2223
rect 6660 2217 6780 2223
rect 6932 2217 7292 2223
rect 7300 2217 7356 2223
rect 3272 2214 3320 2216
rect 3272 2206 3276 2214
rect 3286 2206 3292 2214
rect 3300 2206 3306 2214
rect 3316 2206 3320 2214
rect 3272 2204 3320 2206
rect 6344 2214 6392 2216
rect 6344 2206 6348 2214
rect 6358 2206 6364 2214
rect 6372 2206 6378 2214
rect 6388 2206 6392 2214
rect 6344 2204 6392 2206
rect 84 2197 156 2203
rect 244 2197 284 2203
rect 372 2197 396 2203
rect 404 2197 620 2203
rect 628 2197 748 2203
rect 1428 2197 1676 2203
rect 2628 2197 2652 2203
rect 2692 2197 2860 2203
rect 3341 2197 3932 2203
rect 1332 2177 2172 2183
rect 2436 2177 2684 2183
rect 2788 2177 2844 2183
rect 2852 2177 3164 2183
rect 3341 2183 3347 2197
rect 4484 2197 4588 2203
rect 4724 2197 4972 2203
rect 5268 2197 5484 2203
rect 6532 2197 6700 2203
rect 7284 2197 7308 2203
rect 3172 2177 3347 2183
rect 4500 2177 4700 2183
rect 4708 2177 5116 2183
rect 5348 2177 5516 2183
rect 5524 2177 5612 2183
rect 6180 2177 6332 2183
rect 6541 2177 6684 2183
rect 6541 2164 6547 2177
rect 6708 2177 6844 2183
rect 7124 2177 7187 2183
rect 7181 2164 7187 2177
rect 7220 2177 7276 2183
rect 7300 2177 7388 2183
rect 196 2157 492 2163
rect 500 2157 716 2163
rect 724 2157 732 2163
rect 1156 2157 1180 2163
rect 1188 2157 1292 2163
rect 1620 2157 1660 2163
rect 1668 2157 1788 2163
rect 1796 2157 1852 2163
rect 2116 2157 2156 2163
rect 2180 2157 2716 2163
rect 2740 2157 2764 2163
rect 2996 2157 3036 2163
rect 3044 2157 3068 2163
rect 3700 2157 3788 2163
rect 3844 2157 4044 2163
rect 4068 2157 4172 2163
rect 4452 2157 4476 2163
rect 4484 2157 4668 2163
rect 4804 2157 5100 2163
rect 5108 2157 5308 2163
rect 5396 2157 5532 2163
rect 5652 2157 5692 2163
rect 5700 2157 5788 2163
rect 5860 2157 6028 2163
rect 6052 2157 6076 2163
rect 6244 2157 6284 2163
rect 6292 2157 6300 2163
rect 6484 2157 6540 2163
rect 6580 2157 6732 2163
rect 6756 2157 6796 2163
rect 7076 2157 7155 2163
rect 7149 2144 7155 2157
rect 7188 2157 7372 2163
rect 7380 2157 7468 2163
rect 132 2137 204 2143
rect 228 2137 524 2143
rect 644 2137 732 2143
rect 996 2137 1148 2143
rect 1156 2137 1244 2143
rect 1284 2137 1308 2143
rect 1588 2137 1708 2143
rect 2116 2137 2188 2143
rect 2196 2137 2380 2143
rect 2564 2137 2748 2143
rect 2772 2137 2924 2143
rect 2932 2137 2972 2143
rect 3684 2137 4124 2143
rect 4132 2137 4188 2143
rect 4244 2137 4284 2143
rect 4324 2137 4412 2143
rect 4996 2137 5036 2143
rect 5044 2137 5100 2143
rect 5108 2137 5180 2143
rect 5476 2137 5548 2143
rect 6084 2137 6204 2143
rect 6228 2137 6236 2143
rect 6372 2137 6700 2143
rect 6788 2137 6860 2143
rect 7012 2137 7132 2143
rect 7156 2137 7324 2143
rect 7332 2137 7420 2143
rect 7428 2137 7500 2143
rect 7556 2137 7740 2143
rect 7748 2137 7948 2143
rect 116 2117 140 2123
rect 180 2117 252 2123
rect 308 2117 460 2123
rect 580 2117 668 2123
rect 692 2117 812 2123
rect 1028 2117 1212 2123
rect 1684 2117 1820 2123
rect 1860 2117 1932 2123
rect 2180 2117 2316 2123
rect 2596 2117 2748 2123
rect 2756 2117 2892 2123
rect 2900 2117 3020 2123
rect 3316 2117 3468 2123
rect 3604 2117 3660 2123
rect 3828 2117 3948 2123
rect 3956 2117 4092 2123
rect 4388 2117 4668 2123
rect 4964 2117 5068 2123
rect 5284 2117 5372 2123
rect 5572 2117 5676 2123
rect 5732 2117 5820 2123
rect 6452 2117 6892 2123
rect 6916 2117 7052 2123
rect 7252 2117 7500 2123
rect 7716 2117 7788 2123
rect 7844 2117 7852 2123
rect 7860 2117 7868 2123
rect 212 2097 348 2103
rect 1812 2097 1884 2103
rect 1892 2097 1948 2103
rect 2692 2097 2764 2103
rect 2788 2097 2812 2103
rect 3172 2097 3420 2103
rect 3428 2097 3500 2103
rect 3636 2097 3836 2103
rect 3844 2097 3900 2103
rect 3908 2097 4028 2103
rect 4036 2097 4060 2103
rect 5668 2097 5900 2103
rect 6324 2097 6444 2103
rect 6452 2097 6524 2103
rect 6724 2097 6748 2103
rect 6852 2097 6908 2103
rect 6916 2097 6956 2103
rect 7044 2097 7228 2103
rect 7236 2097 7356 2103
rect 7716 2097 7772 2103
rect 7812 2097 7836 2103
rect 7876 2097 8060 2103
rect 8164 2097 8195 2103
rect 20 2077 76 2083
rect 84 2077 252 2083
rect 260 2077 284 2083
rect 292 2077 620 2083
rect 628 2077 668 2083
rect 948 2077 1068 2083
rect 1076 2077 1388 2083
rect 1556 2077 1868 2083
rect 2580 2077 2716 2083
rect 2788 2077 2860 2083
rect 2868 2077 2940 2083
rect 2948 2077 3148 2083
rect 3364 2077 3532 2083
rect 3540 2077 3852 2083
rect 4964 2077 5020 2083
rect 5060 2077 5180 2083
rect 5796 2077 5868 2083
rect 5876 2077 6108 2083
rect 6116 2077 6716 2083
rect 6772 2077 6876 2083
rect 7156 2077 7772 2083
rect 7812 2077 7932 2083
rect 1300 2057 2812 2063
rect 3988 2057 3996 2063
rect 4004 2057 4236 2063
rect 6484 2057 6668 2063
rect 6676 2057 6812 2063
rect 1348 2037 1820 2043
rect 3988 2037 5436 2043
rect 5444 2037 5580 2043
rect 5588 2037 5916 2043
rect 6644 2037 6668 2043
rect 2308 2017 3276 2023
rect 3284 2017 3452 2023
rect 3668 2017 3756 2023
rect 3972 2017 4540 2023
rect 6260 2017 6924 2023
rect 1736 2014 1784 2016
rect 1736 2006 1740 2014
rect 1750 2006 1756 2014
rect 1764 2006 1770 2014
rect 1780 2006 1784 2014
rect 1736 2004 1784 2006
rect 4808 2014 4856 2016
rect 4808 2006 4812 2014
rect 4822 2006 4828 2014
rect 4836 2006 4842 2014
rect 4852 2006 4856 2014
rect 4808 2004 4856 2006
rect 1364 1997 1372 2003
rect 2708 1997 2764 2003
rect 3108 1997 3196 2003
rect 3652 1997 3756 2003
rect 3940 1997 4156 2003
rect 5316 1997 5756 2003
rect 6596 1997 6876 2003
rect 7076 1997 7804 2003
rect 916 1977 1228 1983
rect 1316 1977 2828 1983
rect 2836 1977 2876 1983
rect 4148 1977 4284 1983
rect 5444 1977 7276 1983
rect 7332 1977 7964 1983
rect 660 1957 844 1963
rect 1412 1957 1452 1963
rect 1460 1957 1596 1963
rect 2276 1957 2332 1963
rect 2500 1957 2556 1963
rect 2564 1957 2796 1963
rect 2804 1957 2844 1963
rect 2852 1957 3356 1963
rect 3396 1957 3468 1963
rect 3476 1957 3708 1963
rect 3764 1957 3820 1963
rect 3908 1957 3948 1963
rect 4084 1957 5948 1963
rect 5956 1957 6076 1963
rect 7316 1957 7452 1963
rect 356 1937 636 1943
rect 676 1937 716 1943
rect 1028 1937 1235 1943
rect 212 1917 220 1923
rect 804 1917 844 1923
rect 852 1917 908 1923
rect 916 1917 1004 1923
rect 1012 1917 1084 1923
rect 1172 1917 1212 1923
rect 1229 1923 1235 1937
rect 1252 1937 1596 1943
rect 2148 1937 2316 1943
rect 2324 1937 2444 1943
rect 3108 1937 3228 1943
rect 3732 1937 4012 1943
rect 4020 1937 4316 1943
rect 4724 1937 4876 1943
rect 4900 1937 5052 1943
rect 5060 1937 5324 1943
rect 6276 1937 6556 1943
rect 7732 1937 8076 1943
rect 8164 1937 8195 1943
rect 1229 1917 1244 1923
rect 1332 1917 1372 1923
rect 1380 1917 1468 1923
rect 2228 1917 2396 1923
rect 3076 1917 3132 1923
rect 3268 1917 3340 1923
rect 3796 1917 3868 1923
rect 4004 1917 4044 1923
rect 4109 1917 4188 1923
rect 4109 1904 4115 1917
rect 4516 1917 4588 1923
rect 5124 1917 5148 1923
rect 5396 1917 5468 1923
rect 5508 1917 5660 1923
rect 5700 1917 5836 1923
rect 6292 1917 6412 1923
rect 6788 1917 6844 1923
rect 6852 1917 6924 1923
rect 7028 1917 7324 1923
rect 7460 1917 7500 1923
rect 7844 1917 7868 1923
rect 7956 1917 8051 1923
rect 36 1897 60 1903
rect 388 1897 428 1903
rect 676 1897 764 1903
rect 772 1897 892 1903
rect 916 1897 972 1903
rect 980 1897 1068 1903
rect 1076 1897 1116 1903
rect 1188 1897 1372 1903
rect 1748 1897 1788 1903
rect 1956 1897 2204 1903
rect 2404 1897 2524 1903
rect 2980 1897 3036 1903
rect 3092 1897 3180 1903
rect 3188 1897 3596 1903
rect 3620 1897 3692 1903
rect 3796 1897 3836 1903
rect 3844 1897 4028 1903
rect 4036 1897 4108 1903
rect 4180 1897 4220 1903
rect 4228 1897 4396 1903
rect 4404 1897 4412 1903
rect 4420 1897 4604 1903
rect 4788 1897 4812 1903
rect 4868 1897 4956 1903
rect 5012 1897 5084 1903
rect 5140 1897 5228 1903
rect 5236 1897 5276 1903
rect 5284 1897 5420 1903
rect 5476 1897 5500 1903
rect 5556 1897 5564 1903
rect 5572 1897 5580 1903
rect 5860 1897 6028 1903
rect 6180 1897 6332 1903
rect 6420 1897 6492 1903
rect 6532 1897 6764 1903
rect 6772 1897 6844 1903
rect 6900 1897 6988 1903
rect 7284 1897 7420 1903
rect 7460 1897 7484 1903
rect 7540 1897 7740 1903
rect 7780 1897 7852 1903
rect 7860 1897 8012 1903
rect 8045 1903 8051 1917
rect 8068 1917 8140 1923
rect 8045 1897 8195 1903
rect 372 1877 492 1883
rect 1044 1877 1196 1883
rect 1364 1877 1436 1883
rect 1684 1877 1772 1883
rect 1940 1877 2044 1883
rect 2196 1877 2332 1883
rect 2340 1877 2380 1883
rect 2388 1877 2524 1883
rect 2532 1877 2572 1883
rect 2580 1877 2668 1883
rect 2692 1877 2748 1883
rect 2820 1877 2908 1883
rect 3140 1877 3196 1883
rect 3268 1877 3436 1883
rect 3844 1877 3884 1883
rect 3924 1877 3964 1883
rect 4116 1877 5340 1883
rect 5428 1877 5564 1883
rect 5652 1877 5708 1883
rect 6532 1877 6572 1883
rect 6724 1877 6844 1883
rect 7028 1877 7148 1883
rect 7204 1877 7324 1883
rect 7524 1877 7596 1883
rect 7828 1877 7852 1883
rect 7860 1877 8012 1883
rect 100 1857 300 1863
rect 308 1857 460 1863
rect 1300 1857 1356 1863
rect 1364 1857 1484 1863
rect 2196 1857 2588 1863
rect 2596 1857 2652 1863
rect 2708 1857 2812 1863
rect 3012 1857 3180 1863
rect 3188 1857 3388 1863
rect 3396 1857 3820 1863
rect 4068 1857 4364 1863
rect 4500 1857 4620 1863
rect 4820 1857 5372 1863
rect 5524 1857 5628 1863
rect 5636 1857 5724 1863
rect 6452 1857 6588 1863
rect 6612 1857 6796 1863
rect 6884 1857 6988 1863
rect 8004 1857 8044 1863
rect 868 1837 908 1843
rect 916 1837 988 1843
rect 996 1837 1084 1843
rect 1428 1837 1836 1843
rect 2068 1837 2124 1843
rect 2701 1843 2707 1856
rect 2132 1837 2707 1843
rect 2788 1837 2876 1843
rect 2916 1837 3052 1843
rect 3220 1837 3372 1843
rect 3924 1837 4524 1843
rect 4564 1837 4764 1843
rect 4788 1837 5196 1843
rect 5204 1837 5244 1843
rect 5268 1837 5724 1843
rect 5988 1837 6092 1843
rect 6132 1837 6252 1843
rect 6468 1837 6636 1843
rect 6740 1837 7116 1843
rect 900 1817 940 1823
rect 2244 1817 2604 1823
rect 2900 1817 3244 1823
rect 3364 1817 3996 1823
rect 4004 1817 4076 1823
rect 4548 1817 4684 1823
rect 4996 1817 5036 1823
rect 5220 1817 5340 1823
rect 5348 1817 5452 1823
rect 5460 1817 5532 1823
rect 5597 1817 5692 1823
rect 3272 1814 3320 1816
rect 3272 1806 3276 1814
rect 3286 1806 3292 1814
rect 3300 1806 3306 1814
rect 3316 1806 3320 1814
rect 3272 1804 3320 1806
rect 596 1797 636 1803
rect 1844 1797 2060 1803
rect 2548 1797 2828 1803
rect 2836 1797 2940 1803
rect 3460 1797 3644 1803
rect 3652 1797 3740 1803
rect 3780 1797 3852 1803
rect 3860 1797 3932 1803
rect 3940 1797 4060 1803
rect 4276 1797 4396 1803
rect 4452 1797 4476 1803
rect 4612 1797 4652 1803
rect 5060 1797 5116 1803
rect 5124 1797 5260 1803
rect 5332 1797 5356 1803
rect 5597 1803 5603 1817
rect 6344 1814 6392 1816
rect 6344 1806 6348 1814
rect 6358 1806 6364 1814
rect 6372 1806 6378 1814
rect 6388 1806 6392 1814
rect 6344 1804 6392 1806
rect 5476 1797 5603 1803
rect 5620 1797 5660 1803
rect 6820 1797 6892 1803
rect 6900 1797 7260 1803
rect 436 1777 524 1783
rect 532 1777 620 1783
rect 724 1777 828 1783
rect 1188 1777 1308 1783
rect 1876 1777 2108 1783
rect 2436 1777 2492 1783
rect 2516 1777 2588 1783
rect 2596 1777 2876 1783
rect 2884 1777 3068 1783
rect 3252 1777 3324 1783
rect 3444 1777 3628 1783
rect 3636 1777 3763 1783
rect 3757 1764 3763 1777
rect 3780 1777 4124 1783
rect 4260 1777 4339 1783
rect 244 1757 332 1763
rect 340 1757 540 1763
rect 644 1757 732 1763
rect 788 1757 908 1763
rect 932 1757 1052 1763
rect 1380 1757 1436 1763
rect 1668 1757 1692 1763
rect 1844 1757 1964 1763
rect 2276 1757 2396 1763
rect 2724 1757 2844 1763
rect 2884 1757 3036 1763
rect 3060 1757 3196 1763
rect 3284 1757 3356 1763
rect 3380 1757 3500 1763
rect 3508 1757 3660 1763
rect 3764 1757 3804 1763
rect 4125 1763 4131 1776
rect 3828 1757 3907 1763
rect 4125 1757 4316 1763
rect 3901 1744 3907 1757
rect 4333 1763 4339 1777
rect 4356 1777 5004 1783
rect 5028 1777 5084 1783
rect 5412 1777 5708 1783
rect 5716 1777 5948 1783
rect 6148 1777 6444 1783
rect 6580 1777 6684 1783
rect 6708 1777 6892 1783
rect 7220 1777 7404 1783
rect 7412 1777 7564 1783
rect 7924 1777 7948 1783
rect 4333 1757 4380 1763
rect 4468 1757 4476 1763
rect 4644 1757 4700 1763
rect 4996 1757 5068 1763
rect 5236 1757 5324 1763
rect 5636 1757 5756 1763
rect 5892 1757 5932 1763
rect 5940 1757 6012 1763
rect 6404 1757 6476 1763
rect 6484 1757 6540 1763
rect 6596 1757 6620 1763
rect 6740 1757 6828 1763
rect 7124 1757 7180 1763
rect 7380 1757 7516 1763
rect 7988 1757 8012 1763
rect 708 1737 796 1743
rect 804 1737 940 1743
rect 964 1737 1068 1743
rect 1236 1737 1532 1743
rect 1700 1737 1820 1743
rect 2052 1737 2092 1743
rect 2212 1737 2636 1743
rect 2660 1737 2700 1743
rect 2852 1737 2924 1743
rect 3156 1737 3180 1743
rect 3220 1737 3260 1743
rect 3364 1737 3404 1743
rect 3540 1737 3580 1743
rect 3604 1737 3676 1743
rect 3684 1737 3852 1743
rect 3908 1737 4108 1743
rect 4148 1737 4364 1743
rect 5092 1737 5196 1743
rect 5316 1737 5340 1743
rect 5444 1737 5788 1743
rect 6244 1737 6364 1743
rect 6372 1737 6492 1743
rect 6500 1737 6508 1743
rect 6516 1737 6604 1743
rect 6612 1737 6668 1743
rect 7892 1737 7980 1743
rect 340 1717 444 1723
rect 772 1717 796 1723
rect 900 1717 1004 1723
rect 1268 1717 1324 1723
rect 1732 1717 1900 1723
rect 2036 1717 2076 1723
rect 2820 1717 3100 1723
rect 3108 1717 4028 1723
rect 4100 1717 4444 1723
rect 4628 1717 4668 1723
rect 4676 1717 4716 1723
rect 5044 1717 5244 1723
rect 5268 1717 5596 1723
rect 5700 1717 5820 1723
rect 6452 1717 6524 1723
rect 6532 1717 6748 1723
rect 6980 1717 7084 1723
rect 7348 1717 7436 1723
rect 68 1697 172 1703
rect 692 1697 956 1703
rect 1124 1697 1324 1703
rect 1460 1697 1708 1703
rect 2084 1697 2188 1703
rect 2340 1697 2716 1703
rect 2740 1697 3148 1703
rect 3172 1697 3212 1703
rect 3268 1697 3772 1703
rect 3796 1697 3820 1703
rect 4429 1697 4492 1703
rect 36 1677 124 1683
rect 548 1677 604 1683
rect 1060 1677 1388 1683
rect 1604 1677 1644 1683
rect 2100 1677 2156 1683
rect 2164 1677 2204 1683
rect 2452 1677 2604 1683
rect 2612 1677 2668 1683
rect 2676 1677 2892 1683
rect 2900 1677 2956 1683
rect 3028 1677 3420 1683
rect 3428 1677 3500 1683
rect 3789 1683 3795 1696
rect 3508 1677 3795 1683
rect 4020 1677 4188 1683
rect 4429 1683 4435 1697
rect 4516 1697 6476 1703
rect 6500 1697 6588 1703
rect 6868 1697 6972 1703
rect 7316 1697 7356 1703
rect 4196 1677 4435 1683
rect 4452 1677 4828 1683
rect 4932 1677 5404 1683
rect 6180 1677 6636 1683
rect 6644 1677 6700 1683
rect 6884 1677 7228 1683
rect 7236 1677 7436 1683
rect 1332 1657 1500 1663
rect 2548 1657 2684 1663
rect 3028 1657 3404 1663
rect 3412 1657 3740 1663
rect 3748 1657 3868 1663
rect 3876 1657 3948 1663
rect 4388 1657 4412 1663
rect 6340 1657 6428 1663
rect 6596 1657 6652 1663
rect 6660 1657 6780 1663
rect 7220 1657 7580 1663
rect 436 1637 460 1643
rect 1476 1637 1500 1643
rect 2020 1637 2348 1643
rect 2356 1637 2460 1643
rect 2532 1637 2684 1643
rect 2788 1637 2988 1643
rect 2996 1637 3116 1643
rect 3220 1637 3452 1643
rect 3460 1637 3516 1643
rect 3588 1637 3932 1643
rect 4084 1637 6876 1643
rect 7156 1637 7180 1643
rect 7412 1637 7644 1643
rect 708 1617 1676 1623
rect 2756 1617 3132 1623
rect 3684 1617 4508 1623
rect 6276 1617 6620 1623
rect 1736 1614 1784 1616
rect 1736 1606 1740 1614
rect 1750 1606 1756 1614
rect 1764 1606 1770 1614
rect 1780 1606 1784 1614
rect 1736 1604 1784 1606
rect 4808 1614 4856 1616
rect 4808 1606 4812 1614
rect 4822 1606 4828 1614
rect 4836 1606 4842 1614
rect 4852 1606 4856 1614
rect 4808 1604 4856 1606
rect 916 1597 1548 1603
rect 2868 1597 3564 1603
rect 3716 1597 4076 1603
rect 4100 1597 4412 1603
rect 6164 1597 6460 1603
rect 6484 1597 7196 1603
rect 1076 1577 1164 1583
rect 1693 1577 1836 1583
rect 1693 1564 1699 1577
rect 2596 1577 2764 1583
rect 3012 1577 4579 1583
rect 228 1557 284 1563
rect 292 1557 396 1563
rect 1108 1557 1340 1563
rect 1549 1557 1692 1563
rect 1549 1544 1555 1557
rect 1716 1557 1948 1563
rect 3604 1557 3980 1563
rect 4052 1557 4252 1563
rect 4573 1563 4579 1577
rect 4660 1577 4988 1583
rect 5044 1577 5084 1583
rect 5268 1577 5692 1583
rect 6436 1577 6732 1583
rect 7012 1577 7052 1583
rect 7060 1577 7100 1583
rect 4573 1557 5276 1563
rect 5412 1557 5708 1563
rect 6116 1557 6396 1563
rect 6948 1557 7084 1563
rect 100 1537 316 1543
rect 1140 1537 1228 1543
rect 1348 1537 1548 1543
rect 1588 1537 1868 1543
rect 1876 1537 1916 1543
rect 3268 1537 3724 1543
rect 3940 1537 4204 1543
rect 4708 1537 4892 1543
rect 5700 1537 5980 1543
rect 6132 1537 6252 1543
rect 6532 1537 6540 1543
rect 6868 1537 6988 1543
rect 7732 1537 7772 1543
rect 7812 1537 7900 1543
rect 148 1517 236 1523
rect 244 1517 412 1523
rect 1028 1517 1164 1523
rect 1229 1523 1235 1536
rect 1229 1517 1468 1523
rect 1684 1517 1708 1523
rect 1764 1517 1804 1523
rect 2292 1517 2300 1523
rect 2676 1517 3004 1523
rect 3236 1517 3532 1523
rect 4052 1517 4140 1523
rect 4180 1517 4316 1523
rect 4324 1517 4428 1523
rect 4596 1517 4748 1523
rect 5124 1517 5228 1523
rect 5556 1517 6707 1523
rect 164 1497 220 1503
rect 340 1497 492 1503
rect 532 1497 572 1503
rect 740 1497 764 1503
rect 836 1497 972 1503
rect 1060 1497 1148 1503
rect 1204 1497 1228 1503
rect 1268 1497 1404 1503
rect 1444 1497 1516 1503
rect 1524 1497 1564 1503
rect 1572 1497 1772 1503
rect 1780 1497 1884 1503
rect 2052 1497 2076 1503
rect 2180 1497 2284 1503
rect 2292 1497 2316 1503
rect 2836 1497 3068 1503
rect 3108 1497 3356 1503
rect 3460 1497 3468 1503
rect 3476 1497 3852 1503
rect 3860 1497 3964 1503
rect 4164 1497 4284 1503
rect 4292 1497 4364 1503
rect 4372 1497 4380 1503
rect 4388 1497 4396 1503
rect 4500 1497 4524 1503
rect 4708 1497 4716 1503
rect 4724 1497 4732 1503
rect 4900 1497 4940 1503
rect 5236 1497 5292 1503
rect 5636 1497 5756 1503
rect 5780 1497 5804 1503
rect 6228 1497 6300 1503
rect 6420 1497 6428 1503
rect 6516 1497 6572 1503
rect 6701 1503 6707 1517
rect 6724 1517 6748 1523
rect 6756 1517 6780 1523
rect 6845 1517 7500 1523
rect 6845 1503 6851 1517
rect 7508 1517 7548 1523
rect 7636 1517 7692 1523
rect 7700 1517 7820 1523
rect 7876 1517 7932 1523
rect 7940 1517 7964 1523
rect 6701 1497 6851 1503
rect 6868 1497 6972 1503
rect 7092 1497 7196 1503
rect 7268 1497 7484 1503
rect 7588 1497 7996 1503
rect 8004 1497 8108 1503
rect 20 1477 76 1483
rect 116 1477 156 1483
rect 164 1477 268 1483
rect 356 1477 380 1483
rect 420 1477 540 1483
rect 692 1477 700 1483
rect 1156 1477 1212 1483
rect 1236 1477 1356 1483
rect 1492 1477 1708 1483
rect 1716 1477 1820 1483
rect 2308 1477 2556 1483
rect 2724 1477 2860 1483
rect 2868 1477 3052 1483
rect 3252 1477 3420 1483
rect 3636 1477 3692 1483
rect 3924 1477 4188 1483
rect 4212 1477 4316 1483
rect 4372 1477 4396 1483
rect 4404 1477 4444 1483
rect 4724 1477 4764 1483
rect 4772 1477 4876 1483
rect 4884 1477 4972 1483
rect 5108 1477 5340 1483
rect 5604 1477 5820 1483
rect 5828 1477 5884 1483
rect 5940 1477 6284 1483
rect 6548 1477 6652 1483
rect 6788 1477 6828 1483
rect 6836 1477 6876 1483
rect 6980 1477 7292 1483
rect 7300 1477 7420 1483
rect 7476 1477 7596 1483
rect 7604 1477 7660 1483
rect 7668 1477 7740 1483
rect 7748 1477 7852 1483
rect 7860 1477 7884 1483
rect 7892 1477 8012 1483
rect 36 1457 124 1463
rect 532 1457 556 1463
rect 1172 1457 1340 1463
rect 1348 1457 1420 1463
rect 1428 1457 1580 1463
rect 1604 1457 1900 1463
rect 1908 1457 1948 1463
rect 3604 1457 3884 1463
rect 3988 1457 4060 1463
rect 4084 1457 4108 1463
rect 4436 1457 4620 1463
rect 4996 1457 5180 1463
rect 6132 1457 6188 1463
rect 6212 1457 6236 1463
rect 6244 1457 6620 1463
rect 6628 1457 6748 1463
rect 6820 1457 6908 1463
rect 7364 1457 7580 1463
rect 7588 1457 7724 1463
rect 7764 1457 7804 1463
rect 7812 1457 7964 1463
rect 7972 1457 8044 1463
rect 484 1437 556 1443
rect 1284 1437 1308 1443
rect 1316 1437 1500 1443
rect 1540 1437 2268 1443
rect 3364 1437 3548 1443
rect 3556 1437 5484 1443
rect 5860 1437 6684 1443
rect 7684 1437 7772 1443
rect 7908 1437 7932 1443
rect 7940 1437 7948 1443
rect 1716 1417 2124 1423
rect 2260 1417 2300 1423
rect 3844 1417 4076 1423
rect 4116 1417 4300 1423
rect 4308 1417 4460 1423
rect 4548 1417 4604 1423
rect 4612 1417 4812 1423
rect 4820 1417 5020 1423
rect 5348 1417 5500 1423
rect 5508 1417 5772 1423
rect 5780 1417 5948 1423
rect 6580 1417 6748 1423
rect 6980 1417 7196 1423
rect 7716 1417 7756 1423
rect 3272 1414 3320 1416
rect 3272 1406 3276 1414
rect 3286 1406 3292 1414
rect 3300 1406 3306 1414
rect 3316 1406 3320 1414
rect 3272 1404 3320 1406
rect 6344 1414 6392 1416
rect 6344 1406 6348 1414
rect 6358 1406 6364 1414
rect 6372 1406 6378 1414
rect 6388 1406 6392 1414
rect 6344 1404 6392 1406
rect 900 1397 924 1403
rect 932 1397 1148 1403
rect 1348 1397 1484 1403
rect 2068 1397 2172 1403
rect 3812 1397 4204 1403
rect 4436 1397 4492 1403
rect 4676 1397 4732 1403
rect 5444 1397 5532 1403
rect 5540 1397 5580 1403
rect 5588 1397 5628 1403
rect 5636 1397 5900 1403
rect 5908 1397 5964 1403
rect 5972 1397 6108 1403
rect 6676 1397 7052 1403
rect 7076 1397 7116 1403
rect 7124 1397 7308 1403
rect 548 1377 684 1383
rect 1188 1377 1292 1383
rect 1300 1377 1468 1383
rect 1476 1377 1612 1383
rect 1620 1377 1692 1383
rect 1972 1377 2028 1383
rect 2333 1377 2492 1383
rect 2333 1364 2339 1377
rect 3396 1377 3596 1383
rect 3732 1377 3820 1383
rect 3828 1377 3923 1383
rect 132 1357 380 1363
rect 404 1357 460 1363
rect 1028 1357 1100 1363
rect 1108 1357 1164 1363
rect 1332 1357 2220 1363
rect 2228 1357 2252 1363
rect 2260 1357 2332 1363
rect 2436 1357 2876 1363
rect 2884 1357 2908 1363
rect 3540 1357 3868 1363
rect 3876 1357 3900 1363
rect 3917 1363 3923 1377
rect 4084 1377 4348 1383
rect 4724 1377 4780 1383
rect 5396 1377 5452 1383
rect 5492 1377 5580 1383
rect 5588 1377 5756 1383
rect 5764 1377 5788 1383
rect 6292 1377 6460 1383
rect 6468 1377 6556 1383
rect 7540 1377 8028 1383
rect 3917 1357 5244 1363
rect 5261 1357 5276 1363
rect 20 1337 412 1343
rect 420 1337 572 1343
rect 580 1337 588 1343
rect 596 1337 636 1343
rect 1140 1337 1196 1343
rect 1204 1337 1340 1343
rect 1492 1337 1596 1343
rect 2132 1337 2188 1343
rect 2900 1337 3100 1343
rect 3460 1337 3516 1343
rect 4020 1337 4124 1343
rect 4173 1337 4348 1343
rect 4173 1324 4179 1337
rect 4916 1337 4940 1343
rect 5261 1343 5267 1357
rect 5492 1357 5660 1363
rect 5748 1357 5868 1363
rect 5892 1357 5916 1363
rect 5924 1357 6044 1363
rect 6132 1357 6444 1363
rect 6452 1357 6460 1363
rect 6468 1357 6588 1363
rect 7828 1357 7900 1363
rect 5204 1337 5267 1343
rect 5284 1337 5308 1343
rect 5316 1337 5468 1343
rect 5476 1337 5516 1343
rect 5524 1337 5548 1343
rect 6164 1337 6236 1343
rect 6692 1337 6908 1343
rect 7412 1337 7532 1343
rect 7956 1337 8044 1343
rect 52 1317 140 1323
rect 180 1317 236 1323
rect 388 1317 428 1323
rect 468 1317 492 1323
rect 580 1317 796 1323
rect 804 1317 876 1323
rect 1380 1317 1612 1323
rect 1860 1317 1916 1323
rect 1956 1317 2076 1323
rect 2340 1317 2412 1323
rect 2420 1317 2492 1323
rect 3044 1317 3132 1323
rect 3236 1317 3356 1323
rect 3636 1317 3740 1323
rect 3972 1317 4060 1323
rect 4068 1317 4172 1323
rect 4196 1317 4332 1323
rect 4340 1317 4364 1323
rect 4468 1317 4524 1323
rect 4724 1317 4876 1323
rect 4916 1317 5020 1323
rect 5172 1317 5196 1323
rect 5252 1317 5276 1323
rect 5284 1317 5724 1323
rect 5732 1317 5772 1323
rect 6196 1317 6220 1323
rect 6685 1323 6691 1336
rect 6564 1317 6691 1323
rect 6804 1317 7100 1323
rect 7108 1317 7180 1323
rect 7188 1317 7356 1323
rect 7540 1317 7628 1323
rect 7700 1317 7836 1323
rect 7924 1317 8012 1323
rect 372 1297 444 1303
rect 452 1297 556 1303
rect 564 1297 620 1303
rect 1060 1297 1276 1303
rect 1412 1297 1436 1303
rect 1604 1297 1660 1303
rect 1924 1297 1980 1303
rect 2164 1297 2652 1303
rect 3076 1297 3212 1303
rect 3220 1297 3388 1303
rect 3412 1297 3436 1303
rect 3748 1297 3980 1303
rect 4212 1297 4460 1303
rect 4788 1297 5148 1303
rect 5652 1297 5692 1303
rect 5700 1297 5820 1303
rect 5828 1297 6156 1303
rect 6996 1297 7100 1303
rect 7636 1297 7708 1303
rect 7764 1297 7932 1303
rect 180 1277 300 1283
rect 308 1277 572 1283
rect 1476 1277 1564 1283
rect 1732 1277 1980 1283
rect 1988 1277 2236 1283
rect 2628 1277 2668 1283
rect 3124 1277 3276 1283
rect 3508 1277 3884 1283
rect 3940 1277 4044 1283
rect 4052 1277 4268 1283
rect 4276 1277 4316 1283
rect 4324 1277 4556 1283
rect 4884 1277 4924 1283
rect 4948 1277 5212 1283
rect 6484 1277 6636 1283
rect 6644 1277 6828 1283
rect 6900 1277 6956 1283
rect 7252 1277 7340 1283
rect 7524 1277 7644 1283
rect 7780 1277 7884 1283
rect 7892 1277 7948 1283
rect 276 1257 364 1263
rect 372 1257 492 1263
rect 4244 1257 4284 1263
rect 4388 1257 4492 1263
rect 4868 1257 4988 1263
rect 5444 1257 5676 1263
rect 5684 1257 5868 1263
rect 6596 1257 6620 1263
rect 6628 1257 6924 1263
rect 2356 1237 2572 1243
rect 2644 1237 5324 1243
rect 5332 1237 5612 1243
rect 5620 1237 5708 1243
rect 5716 1237 5756 1243
rect 5764 1237 5836 1243
rect 5844 1237 5948 1243
rect 6356 1237 6428 1243
rect 6436 1237 6620 1243
rect 6676 1237 6700 1243
rect 6708 1237 6812 1243
rect 6820 1237 7084 1243
rect 2228 1217 2579 1223
rect 1736 1214 1784 1216
rect 1736 1206 1740 1214
rect 1750 1206 1756 1214
rect 1764 1206 1770 1214
rect 1780 1206 1784 1214
rect 1736 1204 1784 1206
rect 868 1197 1020 1203
rect 2052 1197 2140 1203
rect 2148 1197 2396 1203
rect 2573 1203 2579 1217
rect 2596 1217 2796 1223
rect 3796 1217 4236 1223
rect 5156 1217 5308 1223
rect 6068 1217 6972 1223
rect 4808 1214 4856 1216
rect 4808 1206 4812 1214
rect 4822 1206 4828 1214
rect 4836 1206 4842 1214
rect 4852 1206 4856 1214
rect 4808 1204 4856 1206
rect 2573 1197 2796 1203
rect 3364 1197 3564 1203
rect 5076 1197 5388 1203
rect 5828 1197 6204 1203
rect 6788 1197 7244 1203
rect 7988 1197 8012 1203
rect 612 1177 1276 1183
rect 1668 1177 2044 1183
rect 2420 1177 2460 1183
rect 2468 1177 2604 1183
rect 3156 1177 3564 1183
rect 3604 1177 3756 1183
rect 4196 1177 4220 1183
rect 4260 1177 5164 1183
rect 5956 1177 6108 1183
rect 6116 1177 6220 1183
rect 6564 1177 6748 1183
rect 372 1157 908 1163
rect 1588 1157 1932 1163
rect 2036 1157 2316 1163
rect 2404 1157 2476 1163
rect 2884 1157 3068 1163
rect 3076 1157 3795 1163
rect 772 1137 860 1143
rect 1028 1137 1100 1143
rect 1108 1137 1276 1143
rect 1284 1137 2124 1143
rect 2340 1137 2364 1143
rect 2372 1137 2508 1143
rect 2628 1137 2684 1143
rect 3412 1137 3548 1143
rect 3700 1137 3772 1143
rect 3789 1143 3795 1157
rect 3892 1157 4092 1163
rect 4756 1157 4796 1163
rect 5348 1157 5404 1163
rect 5524 1157 5900 1163
rect 7716 1157 8060 1163
rect 8068 1157 8140 1163
rect 3789 1137 5628 1143
rect 5636 1137 5980 1143
rect 6324 1137 6604 1143
rect 6772 1137 6860 1143
rect 6932 1137 7212 1143
rect 7524 1137 7596 1143
rect 7604 1137 7612 1143
rect 7652 1137 7980 1143
rect 356 1117 428 1123
rect 676 1117 732 1123
rect 749 1117 908 1123
rect 404 1097 412 1103
rect 749 1103 755 1117
rect 916 1117 988 1123
rect 1556 1117 1756 1123
rect 2324 1117 2412 1123
rect 2436 1117 2828 1123
rect 4020 1117 4044 1123
rect 4660 1117 4732 1123
rect 4772 1117 4956 1123
rect 4996 1117 5052 1123
rect 5172 1117 5244 1123
rect 5252 1117 5372 1123
rect 5716 1117 5788 1123
rect 5876 1117 5916 1123
rect 6084 1117 6236 1123
rect 6276 1117 6476 1123
rect 6516 1117 6652 1123
rect 6804 1117 6956 1123
rect 7188 1117 7244 1123
rect 7444 1117 7660 1123
rect 724 1097 755 1103
rect 868 1097 972 1103
rect 1332 1097 1372 1103
rect 1460 1097 1667 1103
rect 1661 1084 1667 1097
rect 2100 1097 2108 1103
rect 2164 1097 2204 1103
rect 2372 1097 2412 1103
rect 2500 1097 2540 1103
rect 2660 1097 2732 1103
rect 2820 1097 2940 1103
rect 3252 1097 3292 1103
rect 3396 1097 3436 1103
rect 3444 1097 3660 1103
rect 3876 1097 3964 1103
rect 3988 1097 4140 1103
rect 4260 1097 4348 1103
rect 4532 1097 4908 1103
rect 4932 1097 5004 1103
rect 5092 1097 5180 1103
rect 5220 1097 5244 1103
rect 5268 1097 5340 1103
rect 5684 1097 5708 1103
rect 5940 1097 6172 1103
rect 6196 1097 6268 1103
rect 6452 1097 6572 1103
rect 6580 1097 6732 1103
rect 6740 1097 7372 1103
rect 7380 1097 7548 1103
rect 7556 1097 7676 1103
rect 7684 1097 7756 1103
rect 7876 1097 7900 1103
rect 644 1077 652 1083
rect 756 1077 780 1083
rect 804 1077 844 1083
rect 884 1077 940 1083
rect 948 1077 1036 1083
rect 1172 1077 1180 1083
rect 1220 1077 1356 1083
rect 1444 1077 1484 1083
rect 1501 1077 1564 1083
rect 1501 1064 1507 1077
rect 1668 1077 1708 1083
rect 2116 1077 2140 1083
rect 2148 1077 2204 1083
rect 2212 1077 2332 1083
rect 2653 1083 2659 1096
rect 2404 1077 2659 1083
rect 2692 1077 2716 1083
rect 2724 1077 3084 1083
rect 3284 1077 3372 1083
rect 3492 1077 3660 1083
rect 3668 1077 3692 1083
rect 3732 1077 3868 1083
rect 3876 1077 4076 1083
rect 4148 1077 4156 1083
rect 4164 1077 4268 1083
rect 4724 1077 4764 1083
rect 4804 1077 4892 1083
rect 5076 1077 5116 1083
rect 5156 1077 5276 1083
rect 5300 1077 5356 1083
rect 5428 1077 5532 1083
rect 5924 1077 6028 1083
rect 6372 1077 6620 1083
rect 6756 1077 6924 1083
rect 7140 1077 7276 1083
rect 7332 1077 7356 1083
rect 7380 1077 7452 1083
rect 7492 1077 7532 1083
rect 7844 1077 7868 1083
rect 660 1057 1084 1063
rect 1092 1057 1196 1063
rect 1204 1057 1340 1063
rect 1396 1057 1500 1063
rect 1844 1057 2012 1063
rect 2196 1057 2380 1063
rect 2500 1057 2668 1063
rect 2852 1057 2908 1063
rect 3220 1057 3532 1063
rect 3540 1057 3612 1063
rect 3684 1057 3884 1063
rect 3940 1057 4028 1063
rect 4084 1057 4204 1063
rect 4740 1057 4908 1063
rect 4916 1057 4988 1063
rect 4996 1057 5020 1063
rect 5028 1057 5084 1063
rect 5092 1057 5100 1063
rect 5604 1057 5772 1063
rect 5780 1057 6092 1063
rect 6301 1057 6332 1063
rect 212 1037 220 1043
rect 228 1037 316 1043
rect 708 1037 812 1043
rect 1236 1037 1404 1043
rect 1412 1037 1452 1043
rect 2020 1037 2060 1043
rect 2260 1037 2300 1043
rect 2308 1037 2444 1043
rect 2452 1037 2636 1043
rect 2788 1037 2812 1043
rect 2964 1037 3356 1043
rect 3364 1037 3468 1043
rect 3476 1037 3564 1043
rect 3572 1037 3708 1043
rect 3844 1037 4236 1043
rect 4468 1037 4748 1043
rect 5188 1037 5436 1043
rect 6301 1043 6307 1057
rect 7428 1057 7500 1063
rect 7700 1057 7724 1063
rect 7732 1057 7820 1063
rect 7860 1057 7964 1063
rect 7972 1057 8108 1063
rect 5636 1037 6307 1043
rect 6324 1037 6348 1043
rect 6484 1037 6812 1043
rect 6820 1037 6876 1043
rect 6884 1037 7148 1043
rect 7364 1037 7436 1043
rect 516 1017 588 1023
rect 756 1017 764 1023
rect 772 1017 828 1023
rect 836 1017 956 1023
rect 964 1017 988 1023
rect 996 1017 1116 1023
rect 1124 1017 1292 1023
rect 1412 1017 1484 1023
rect 2532 1017 2556 1023
rect 2781 1023 2787 1036
rect 2564 1017 2787 1023
rect 2916 1017 3100 1023
rect 3748 1017 3932 1023
rect 3972 1017 4188 1023
rect 4276 1017 4476 1023
rect 4484 1017 4508 1023
rect 4948 1017 5020 1023
rect 5028 1017 5100 1023
rect 5236 1017 5651 1023
rect 3272 1014 3320 1016
rect 3272 1006 3276 1014
rect 3286 1006 3292 1014
rect 3300 1006 3306 1014
rect 3316 1006 3320 1014
rect 3272 1004 3320 1006
rect 5645 1004 5651 1017
rect 6212 1017 6300 1023
rect 6596 1017 6844 1023
rect 6852 1017 6908 1023
rect 7044 1017 7308 1023
rect 7556 1017 7788 1023
rect 8068 1017 8092 1023
rect 6344 1014 6392 1016
rect 6344 1006 6348 1014
rect 6358 1006 6364 1014
rect 6372 1006 6378 1014
rect 6388 1006 6392 1014
rect 6344 1004 6392 1006
rect 420 997 604 1003
rect 1316 997 1420 1003
rect 1444 997 1468 1003
rect 2228 997 3004 1003
rect 3940 997 4348 1003
rect 4612 997 4700 1003
rect 4708 997 4764 1003
rect 5012 997 5260 1003
rect 5652 997 5724 1003
rect 5732 997 5852 1003
rect 7284 997 7740 1003
rect 116 977 236 983
rect 564 977 668 983
rect 1437 983 1443 996
rect 1268 977 1443 983
rect 1492 977 1708 983
rect 2020 977 2204 983
rect 2724 977 2908 983
rect 3060 977 3116 983
rect 3124 977 3228 983
rect 3236 977 3452 983
rect 3805 977 3932 983
rect 3805 964 3811 977
rect 3940 977 3948 983
rect 3956 977 3980 983
rect 4228 977 4412 983
rect 4484 977 4908 983
rect 4916 977 5068 983
rect 5220 977 5468 983
rect 5476 977 5916 983
rect 6276 977 7132 983
rect 7444 977 7564 983
rect 7572 977 7708 983
rect 7908 977 8108 983
rect 52 957 300 963
rect 308 957 355 963
rect 349 944 355 957
rect 948 957 1020 963
rect 1460 957 1500 963
rect 1508 957 1596 963
rect 2644 957 2700 963
rect 2900 957 2924 963
rect 2932 957 3068 963
rect 3188 957 3228 963
rect 3700 957 3740 963
rect 3748 957 3804 963
rect 4132 957 4268 963
rect 4388 957 4428 963
rect 4468 957 4604 963
rect 4612 957 4780 963
rect 4804 957 5052 963
rect 5060 957 5292 963
rect 5492 957 5708 963
rect 6004 957 6300 963
rect 6365 957 6444 963
rect 148 937 188 943
rect 356 937 364 943
rect 660 937 844 943
rect 852 937 1036 943
rect 1044 937 1244 943
rect 1252 937 1276 943
rect 1284 937 1388 943
rect 1396 937 1420 943
rect 1428 937 1612 943
rect 1636 937 1932 943
rect 2436 937 2716 943
rect 3012 937 3132 943
rect 3140 937 3196 943
rect 3236 937 3676 943
rect 3716 937 3756 943
rect 3796 937 3852 943
rect 3860 937 4140 943
rect 4148 937 4300 943
rect 4596 937 4812 943
rect 4980 937 5084 943
rect 5396 937 5532 943
rect 5540 937 5564 943
rect 5572 937 5692 943
rect 5700 937 5772 943
rect 6068 937 6108 943
rect 6116 937 6124 943
rect 6365 943 6371 957
rect 6900 957 6924 963
rect 6932 957 7196 963
rect 7748 957 8012 963
rect 6157 937 6371 943
rect 6157 924 6163 937
rect 6388 937 6476 943
rect 6660 937 6700 943
rect 6980 937 7372 943
rect 7412 937 7516 943
rect 7652 937 7804 943
rect 36 917 92 923
rect 164 917 204 923
rect 276 917 412 923
rect 788 917 876 923
rect 916 917 1164 923
rect 1236 917 1292 923
rect 1348 917 1379 923
rect 68 897 172 903
rect 212 897 428 903
rect 596 897 684 903
rect 1012 897 1100 903
rect 1188 897 1212 903
rect 1268 897 1356 903
rect 1373 903 1379 917
rect 1396 917 1404 923
rect 1444 917 1660 923
rect 2148 917 2172 923
rect 2692 917 2780 923
rect 2980 917 3244 923
rect 3252 917 3356 923
rect 3364 917 3500 923
rect 3556 917 3596 923
rect 3604 917 3660 923
rect 3924 917 3964 923
rect 4052 917 4156 923
rect 4356 917 4380 923
rect 4516 917 4684 923
rect 4692 917 4972 923
rect 5364 917 5468 923
rect 5684 917 5804 923
rect 5876 917 5996 923
rect 6004 917 6156 923
rect 6180 917 6236 923
rect 6244 917 6284 923
rect 6660 917 6764 923
rect 7076 917 7404 923
rect 7412 917 7484 923
rect 7588 917 7724 923
rect 7860 917 7884 923
rect 1373 897 1548 903
rect 1604 897 1676 903
rect 1684 897 1724 903
rect 1988 897 2124 903
rect 2132 897 2172 903
rect 2692 897 2748 903
rect 3268 897 3436 903
rect 3924 897 4108 903
rect 4564 897 4748 903
rect 4788 897 4924 903
rect 4964 897 5132 903
rect 5668 897 5868 903
rect 6180 897 6284 903
rect 6452 897 6652 903
rect 6660 897 6732 903
rect 7060 897 7308 903
rect 7748 897 7852 903
rect 7892 897 7996 903
rect 20 877 140 883
rect 292 877 316 883
rect 356 877 396 883
rect 644 877 796 883
rect 804 877 860 883
rect 868 877 972 883
rect 1460 877 1644 883
rect 1652 877 1756 883
rect 3844 877 3884 883
rect 3892 877 3900 883
rect 4052 877 4092 883
rect 4212 877 4540 883
rect 4548 877 5212 883
rect 5316 877 5420 883
rect 5748 877 5932 883
rect 5940 877 6140 883
rect 6548 877 6604 883
rect 7348 877 7388 883
rect 7396 877 7468 883
rect 7508 877 7628 883
rect 84 857 364 863
rect 628 857 1228 863
rect 1380 857 2908 863
rect 3076 857 3404 863
rect 3412 857 3644 863
rect 3652 857 3676 863
rect 3876 857 3996 863
rect 4004 857 4028 863
rect 4628 857 4652 863
rect 4660 857 4796 863
rect 4900 857 6940 863
rect 7252 857 7484 863
rect 1716 837 1740 843
rect 2628 837 4844 843
rect 4868 837 4988 843
rect 6941 843 6947 856
rect 6941 837 7372 843
rect 7716 837 7756 843
rect 2068 817 2684 823
rect 3188 817 3372 823
rect 4116 817 4412 823
rect 5524 817 5564 823
rect 5572 817 5612 823
rect 5620 817 5932 823
rect 1736 814 1784 816
rect 1736 806 1740 814
rect 1750 806 1756 814
rect 1764 806 1770 814
rect 1780 806 1784 814
rect 1736 804 1784 806
rect 4808 814 4856 816
rect 4808 806 4812 814
rect 4822 806 4828 814
rect 4836 806 4842 814
rect 4852 806 4856 814
rect 4808 804 4856 806
rect 3972 797 4108 803
rect 4308 797 4540 803
rect 244 777 364 783
rect 372 777 396 783
rect 404 777 588 783
rect 596 777 604 783
rect 3092 777 3132 783
rect 3668 777 4268 783
rect 4484 777 4556 783
rect 132 757 524 763
rect 1508 757 1580 763
rect 2356 757 2492 763
rect 2500 757 2572 763
rect 3796 757 4252 763
rect 5140 757 5196 763
rect 7124 757 7212 763
rect 7220 757 7420 763
rect 36 737 252 743
rect 260 737 284 743
rect 1300 737 2204 743
rect 2212 737 2268 743
rect 2276 737 2540 743
rect 2548 737 2572 743
rect 2580 737 2684 743
rect 2852 737 3004 743
rect 3060 737 3340 743
rect 3716 737 4236 743
rect 5140 737 5228 743
rect 5572 737 6140 743
rect 6436 737 6492 743
rect 6500 737 6748 743
rect 6756 737 7004 743
rect 7012 737 7180 743
rect 8068 737 8076 743
rect 228 717 316 723
rect 468 717 684 723
rect 1348 717 1372 723
rect 1540 717 1644 723
rect 1684 717 1804 723
rect 2228 717 2284 723
rect 2340 717 2380 723
rect 2420 717 2476 723
rect 2612 717 2700 723
rect 2852 717 2924 723
rect 3636 717 3852 723
rect 3860 717 3868 723
rect 3908 717 4156 723
rect 5076 717 5100 723
rect 5188 717 5532 723
rect 5956 717 5980 723
rect 6404 717 6940 723
rect 7380 717 7484 723
rect 7524 717 7596 723
rect 7812 717 7852 723
rect 7860 717 7980 723
rect 8068 717 8108 723
rect 20 697 76 703
rect 84 697 172 703
rect 308 697 332 703
rect 436 697 460 703
rect 916 697 1036 703
rect 1396 697 1436 703
rect 1540 697 1548 703
rect 1636 697 1660 703
rect 1684 697 1772 703
rect 1796 697 1916 703
rect 2285 703 2291 716
rect 2285 697 2428 703
rect 2452 697 2476 703
rect 2596 697 2748 703
rect 2772 697 2828 703
rect 2836 697 2940 703
rect 3348 697 3516 703
rect 3700 697 3708 703
rect 3940 697 4012 703
rect 4036 697 4092 703
rect 4116 697 4140 703
rect 4788 697 4844 703
rect 5076 697 5340 703
rect 5588 697 6012 703
rect 6196 697 6332 703
rect 6340 697 6444 703
rect 6452 697 6524 703
rect 6532 697 6620 703
rect 6660 697 6780 703
rect 6820 697 6876 703
rect 7124 697 7164 703
rect 7172 697 7244 703
rect 7252 697 7420 703
rect 7428 697 7788 703
rect 8020 697 8092 703
rect 180 677 220 683
rect 260 677 348 683
rect 500 677 700 683
rect 1204 677 1228 683
rect 1236 677 1452 683
rect 1460 677 1500 683
rect 2244 677 2268 683
rect 2340 677 2556 683
rect 2564 677 2668 683
rect 2676 677 2780 683
rect 2932 677 3036 683
rect 3268 677 3484 683
rect 3764 677 3804 683
rect 3812 677 4076 683
rect 4084 677 4188 683
rect 4308 677 4380 683
rect 4388 677 4652 683
rect 4692 677 4700 683
rect 4996 677 5148 683
rect 5300 677 5484 683
rect 5492 677 5788 683
rect 6484 677 6732 683
rect 7060 677 7276 683
rect 7332 677 7372 683
rect 7412 677 7452 683
rect 7460 677 7548 683
rect 7780 677 7804 683
rect 7844 677 7868 683
rect 7988 677 8108 683
rect 628 657 812 663
rect 1492 657 1692 663
rect 1860 657 1980 663
rect 2324 657 2716 663
rect 3140 657 3452 663
rect 3716 657 3740 663
rect 3748 657 3820 663
rect 3972 657 4284 663
rect 4292 657 4316 663
rect 4692 657 4876 663
rect 4884 657 5388 663
rect 5444 657 5740 663
rect 5748 657 5772 663
rect 5844 657 5900 663
rect 6084 657 6412 663
rect 7076 657 7132 663
rect 7268 657 7468 663
rect 7732 657 7996 663
rect 8004 657 8028 663
rect 8100 657 8156 663
rect 484 637 508 643
rect 516 637 1260 643
rect 1268 637 1292 643
rect 1300 637 1836 643
rect 2292 637 2844 643
rect 3252 637 3788 643
rect 4980 637 5004 643
rect 5012 637 5468 643
rect 5476 637 5804 643
rect 6068 637 6268 643
rect 6276 637 6316 643
rect 7844 637 7964 643
rect 7972 637 8140 643
rect 1220 617 1596 623
rect 1684 617 2284 623
rect 4036 617 4380 623
rect 4916 617 5084 623
rect 5092 617 5148 623
rect 5812 617 5868 623
rect 6820 617 6860 623
rect 7924 617 8012 623
rect 8020 617 8060 623
rect 3272 614 3320 616
rect 3272 606 3276 614
rect 3286 606 3292 614
rect 3300 606 3306 614
rect 3316 606 3320 614
rect 3272 604 3320 606
rect 6344 614 6392 616
rect 6344 606 6348 614
rect 6358 606 6364 614
rect 6372 606 6378 614
rect 6388 606 6392 614
rect 6344 604 6392 606
rect 20 597 60 603
rect 68 597 380 603
rect 932 597 988 603
rect 996 597 2060 603
rect 2628 597 2668 603
rect 2756 597 2876 603
rect 3652 597 4220 603
rect 5140 597 5564 603
rect 7284 597 7372 603
rect 180 577 396 583
rect 1220 577 1244 583
rect 1412 577 1580 583
rect 2196 577 2412 583
rect 2660 577 3436 583
rect 3652 577 3724 583
rect 3732 577 3932 583
rect 3940 577 4124 583
rect 4253 577 4268 583
rect 4253 564 4259 577
rect 5780 577 5948 583
rect 6292 577 6508 583
rect 6564 577 6684 583
rect 6692 577 6716 583
rect 6724 577 6764 583
rect 6772 577 7020 583
rect 7284 577 7308 583
rect 7492 577 7516 583
rect 292 557 364 563
rect 436 557 636 563
rect 1156 557 1388 563
rect 1572 557 1644 563
rect 2068 557 2124 563
rect 2244 557 2348 563
rect 2452 557 2476 563
rect 2644 557 2748 563
rect 2820 557 3132 563
rect 4324 557 4348 563
rect 4788 557 4924 563
rect 4932 557 4956 563
rect 4964 557 5180 563
rect 5460 557 5564 563
rect 5572 557 5836 563
rect 5940 557 6092 563
rect 6244 557 6316 563
rect 6340 557 6444 563
rect 6452 557 6508 563
rect 6516 557 6540 563
rect 6948 557 7260 563
rect 7268 557 7676 563
rect 148 537 188 543
rect 196 537 204 543
rect 260 537 444 543
rect 1140 537 1532 543
rect 1540 537 1580 543
rect 1876 537 1996 543
rect 2116 537 2268 543
rect 2276 537 2332 543
rect 2340 537 2556 543
rect 2564 537 2652 543
rect 2660 537 2844 543
rect 3348 537 3516 543
rect 3524 537 4028 543
rect 4292 537 4348 543
rect 4900 537 4972 543
rect 4980 537 5004 543
rect 5012 537 5052 543
rect 5060 537 5196 543
rect 5492 537 5628 543
rect 5748 537 5820 543
rect 5828 537 5852 543
rect 5860 537 6012 543
rect 6228 537 6412 543
rect 6532 537 6572 543
rect 6612 537 6812 543
rect 7028 537 7084 543
rect 7444 537 7580 543
rect 356 517 524 523
rect 708 517 780 523
rect 788 517 844 523
rect 1844 517 1980 523
rect 2036 517 2076 523
rect 2260 517 2348 523
rect 2356 517 2604 523
rect 2692 517 2732 523
rect 2740 517 2796 523
rect 2932 517 3084 523
rect 3524 517 3708 523
rect 3876 517 3948 523
rect 4068 517 4188 523
rect 4404 517 4508 523
rect 4772 517 4796 523
rect 4996 517 5100 523
rect 5348 517 5532 523
rect 5684 517 5788 523
rect 6404 517 6588 523
rect 6756 517 6860 523
rect 7044 517 7084 523
rect 7540 517 7628 523
rect 7780 517 7964 523
rect 7988 517 8028 523
rect 8052 517 8060 523
rect 260 497 332 503
rect 340 497 348 503
rect 420 497 492 503
rect 532 497 636 503
rect 820 497 1564 503
rect 1652 497 1676 503
rect 2452 497 2508 503
rect 2580 497 2956 503
rect 3732 497 3852 503
rect 4276 497 4332 503
rect 4404 497 4444 503
rect 5044 497 5260 503
rect 5604 497 5660 503
rect 6125 497 6220 503
rect 6125 484 6131 497
rect 6420 497 6668 503
rect 6676 497 6796 503
rect 7012 497 7180 503
rect 8068 497 8124 503
rect 1652 477 1692 483
rect 1700 477 1932 483
rect 2372 477 2396 483
rect 2404 477 2684 483
rect 3588 477 3804 483
rect 3812 477 4124 483
rect 4180 477 4508 483
rect 5092 477 5244 483
rect 6052 477 6124 483
rect 6164 477 6476 483
rect 6676 477 6716 483
rect 6996 477 7052 483
rect 8036 477 8092 483
rect 420 457 1228 463
rect 1236 457 2028 463
rect 2308 457 3772 463
rect 4212 457 4348 463
rect 4676 457 5100 463
rect 5620 457 5692 463
rect 5700 457 5724 463
rect 5732 457 5916 463
rect 6516 457 6732 463
rect 580 437 764 443
rect 772 437 812 443
rect 2996 437 3260 443
rect 3268 437 3356 443
rect 3444 437 3948 443
rect 4484 437 4556 443
rect 2900 417 3660 423
rect 5428 417 6188 423
rect 1736 414 1784 416
rect 1736 406 1740 414
rect 1750 406 1756 414
rect 1764 406 1770 414
rect 1780 406 1784 414
rect 1736 404 1784 406
rect 4808 414 4856 416
rect 4808 406 4812 414
rect 4822 406 4828 414
rect 4836 406 4842 414
rect 4852 406 4856 414
rect 4808 404 4856 406
rect 3060 397 3756 403
rect 5460 397 6300 403
rect 6308 397 6396 403
rect 7796 397 7852 403
rect 7860 397 7916 403
rect 7924 397 8108 403
rect 2852 377 2908 383
rect 2964 377 3100 383
rect 3124 377 3228 383
rect 3236 377 3644 383
rect 3652 377 3756 383
rect 5204 377 5308 383
rect 6292 377 6444 383
rect 6820 377 7452 383
rect 2596 357 2812 363
rect 2836 357 3020 363
rect 3348 357 3676 363
rect 3812 357 4028 363
rect 4948 357 5020 363
rect 5108 357 5388 363
rect 5396 357 5532 363
rect 5540 357 5980 363
rect 6724 357 6956 363
rect 7028 357 7084 363
rect 7092 357 7132 363
rect 244 337 348 343
rect 372 337 572 343
rect 580 337 620 343
rect 628 337 764 343
rect 1428 337 1564 343
rect 1588 337 1740 343
rect 2452 337 2668 343
rect 2676 337 2908 343
rect 2916 337 2956 343
rect 3364 337 3548 343
rect 3700 337 3916 343
rect 3972 337 4236 343
rect 4580 337 4940 343
rect 5076 337 5116 343
rect 5140 337 5228 343
rect 5668 337 5740 343
rect 6900 337 6924 343
rect 6932 337 7116 343
rect 7124 337 7196 343
rect 260 317 316 323
rect 324 317 444 323
rect 500 317 588 323
rect 1316 317 1452 323
rect 1460 317 1548 323
rect 1684 317 1708 323
rect 1764 317 1932 323
rect 1940 317 2060 323
rect 2388 317 2476 323
rect 2493 317 2716 323
rect 148 297 204 303
rect 356 297 396 303
rect 404 297 444 303
rect 548 297 716 303
rect 884 297 1004 303
rect 1684 297 1820 303
rect 1908 297 2012 303
rect 2020 297 2156 303
rect 2212 297 2396 303
rect 2493 303 2499 317
rect 2756 317 2860 323
rect 3188 317 3292 323
rect 3300 317 3388 323
rect 3492 317 3596 323
rect 3908 317 3932 323
rect 4372 317 4428 323
rect 4468 317 4588 323
rect 4596 317 4620 323
rect 4644 317 4700 323
rect 4996 317 5235 323
rect 5229 304 5235 317
rect 5604 317 5676 323
rect 5780 317 5804 323
rect 5844 317 5900 323
rect 7156 317 7244 323
rect 7508 317 7708 323
rect 7716 317 7884 323
rect 7908 317 7916 323
rect 7924 317 7964 323
rect 2420 297 2499 303
rect 2532 297 2716 303
rect 2724 297 2812 303
rect 2820 297 2988 303
rect 3428 297 3484 303
rect 3556 297 3724 303
rect 3732 297 3884 303
rect 3908 297 4108 303
rect 4436 297 4476 303
rect 4484 297 4604 303
rect 4612 297 4636 303
rect 4660 297 4732 303
rect 5076 297 5164 303
rect 5236 297 5276 303
rect 5476 297 5484 303
rect 5556 297 5628 303
rect 5700 297 5724 303
rect 5732 297 5948 303
rect 6244 297 6460 303
rect 6532 297 6700 303
rect 7140 297 7228 303
rect 7268 297 7324 303
rect 7700 297 7740 303
rect 7812 297 7932 303
rect 7988 297 8060 303
rect 8164 297 8195 303
rect 260 277 396 283
rect 404 277 508 283
rect 516 277 1148 283
rect 1156 277 1244 283
rect 1348 277 1692 283
rect 2548 277 2700 283
rect 2724 277 2828 283
rect 2884 277 3132 283
rect 3412 277 3484 283
rect 3492 277 3532 283
rect 3540 277 3740 283
rect 3748 277 3996 283
rect 4004 277 6012 283
rect 6564 277 6652 283
rect 6660 277 6844 283
rect 6900 277 6972 283
rect 6980 277 7052 283
rect 7428 277 7468 283
rect 7668 277 7708 283
rect 7748 277 7820 283
rect 7828 277 7996 283
rect 8004 277 8028 283
rect 100 257 268 263
rect 324 257 524 263
rect 628 257 652 263
rect 660 257 851 263
rect 845 244 851 257
rect 948 257 1068 263
rect 1172 257 1196 263
rect 1508 257 1628 263
rect 1700 257 1724 263
rect 2484 257 2620 263
rect 2740 257 2764 263
rect 2836 257 3068 263
rect 3636 257 3676 263
rect 3684 257 3708 263
rect 3780 257 3820 263
rect 3892 257 3916 263
rect 3940 257 3980 263
rect 4308 257 4364 263
rect 4500 257 4524 263
rect 4660 257 4684 263
rect 5092 257 5196 263
rect 5204 257 5212 263
rect 5220 257 5292 263
rect 5300 257 5340 263
rect 5636 257 5852 263
rect 6628 257 6796 263
rect 6804 257 6876 263
rect 6884 257 6988 263
rect 6996 257 7036 263
rect 7044 257 7100 263
rect 7972 257 8092 263
rect 852 237 876 243
rect 1540 237 1612 243
rect 1620 237 1884 243
rect 3172 237 3532 243
rect 3540 237 3580 243
rect 3828 237 3868 243
rect 4804 237 4860 243
rect 5620 237 5708 243
rect 5716 237 5788 243
rect 5988 237 6588 243
rect 6596 237 6844 243
rect 6852 237 6860 243
rect 6868 237 7004 243
rect 7620 237 7628 243
rect 7636 237 8012 243
rect 8068 237 8092 243
rect 20 217 188 223
rect 724 217 860 223
rect 1316 217 1388 223
rect 1636 217 1740 223
rect 1748 217 1868 223
rect 3716 217 3836 223
rect 3844 217 3916 223
rect 4356 217 4572 223
rect 4628 217 4876 223
rect 4900 217 5228 223
rect 5236 217 5484 223
rect 6932 217 6956 223
rect 6964 217 7212 223
rect 7860 217 7964 223
rect 3272 214 3320 216
rect 3272 206 3276 214
rect 3286 206 3292 214
rect 3300 206 3306 214
rect 3316 206 3320 214
rect 3272 204 3320 206
rect 6344 214 6392 216
rect 6344 206 6348 214
rect 6358 206 6364 214
rect 6372 206 6378 214
rect 6388 206 6392 214
rect 6344 204 6392 206
rect 404 197 892 203
rect 2244 197 2316 203
rect 2628 197 2803 203
rect 2797 184 2803 197
rect 4308 197 4332 203
rect 4340 197 5724 203
rect 6100 197 6252 203
rect 6724 197 6780 203
rect 6788 197 6988 203
rect 6996 197 7020 203
rect 7876 197 7916 203
rect 596 177 844 183
rect 1517 177 1891 183
rect 1517 164 1523 177
rect 36 157 76 163
rect 148 157 348 163
rect 468 157 716 163
rect 1204 157 1516 163
rect 1540 157 1644 163
rect 1684 157 1708 163
rect 1716 157 1756 163
rect 1885 163 1891 177
rect 1908 177 1996 183
rect 2036 177 2076 183
rect 2116 177 2172 183
rect 2516 177 2556 183
rect 2564 177 2748 183
rect 2804 177 2924 183
rect 2964 177 3004 183
rect 3012 177 3036 183
rect 3396 177 3420 183
rect 3732 177 3740 183
rect 4532 177 4684 183
rect 4724 177 4812 183
rect 4820 177 4924 183
rect 5140 177 5260 183
rect 5268 177 5372 183
rect 5380 177 5468 183
rect 5565 177 5772 183
rect 5565 164 5571 177
rect 6660 177 6732 183
rect 6740 177 6812 183
rect 7764 177 7836 183
rect 7844 177 7996 183
rect 1885 157 1964 163
rect 1972 157 2124 163
rect 2148 157 2172 163
rect 2196 157 2236 163
rect 2644 157 2764 163
rect 2772 157 2892 163
rect 3028 157 3228 163
rect 3780 157 3852 163
rect 4020 157 4060 163
rect 4116 157 4316 163
rect 4516 157 4540 163
rect 4548 157 4588 163
rect 4596 157 4732 163
rect 4852 157 4924 163
rect 5156 157 5187 163
rect 68 137 156 143
rect 164 137 316 143
rect 324 137 588 143
rect 628 137 812 143
rect 836 137 892 143
rect 948 137 1052 143
rect 1620 137 1724 143
rect 1732 137 2156 143
rect 2164 137 2252 143
rect 2260 137 2428 143
rect 2436 137 2524 143
rect 2532 137 2732 143
rect 2756 137 2908 143
rect 2996 137 3132 143
rect 3236 137 3308 143
rect 3444 137 3532 143
rect 3748 137 3788 143
rect 3828 137 4044 143
rect 4084 137 4172 143
rect 4388 137 4428 143
rect 4436 137 4556 143
rect 4580 137 4636 143
rect 4644 137 4764 143
rect 5028 137 5164 143
rect 5181 143 5187 157
rect 5220 157 5308 163
rect 5764 157 5852 163
rect 5940 157 5964 163
rect 5972 157 6108 163
rect 6116 157 6236 163
rect 6292 157 6588 163
rect 6612 157 6668 163
rect 6765 157 6812 163
rect 5181 137 5212 143
rect 5220 137 5260 143
rect 5332 137 5468 143
rect 5588 137 5708 143
rect 5732 137 6476 143
rect 6484 137 6524 143
rect 6548 137 6556 143
rect 6580 137 6636 143
rect 6765 143 6771 157
rect 7284 157 7340 163
rect 7540 157 7852 163
rect 7876 157 7964 163
rect 8020 157 8076 163
rect 6660 137 6771 143
rect 6788 137 6844 143
rect 7124 137 7308 143
rect 7316 137 7404 143
rect 7876 137 7932 143
rect 8068 137 8092 143
rect 84 117 428 123
rect 436 117 476 123
rect 612 117 668 123
rect 740 117 796 123
rect 804 117 956 123
rect 1156 117 1260 123
rect 1332 117 1420 123
rect 1588 117 1692 123
rect 1860 117 1884 123
rect 1892 117 2300 123
rect 2324 117 2780 123
rect 2788 117 2844 123
rect 2916 117 3004 123
rect 3348 117 3452 123
rect 3668 117 3692 123
rect 3700 117 3820 123
rect 3908 117 3948 123
rect 4052 117 5964 123
rect 6404 117 6668 123
rect 6676 117 6764 123
rect 6804 117 6876 123
rect 6900 117 6940 123
rect 6980 117 7052 123
rect 7364 117 7420 123
rect 7604 117 7868 123
rect 7940 117 8060 123
rect 196 97 236 103
rect 244 97 300 103
rect 308 97 412 103
rect 420 97 748 103
rect 884 97 1148 103
rect 1844 97 1900 103
rect 1924 97 1948 103
rect 1956 97 1980 103
rect 2004 97 2044 103
rect 2468 97 2572 103
rect 2612 97 2668 103
rect 3476 97 3692 103
rect 3700 97 3772 103
rect 3876 97 4092 103
rect 4292 97 4396 103
rect 4404 97 4460 103
rect 4468 97 4700 103
rect 4708 97 4748 103
rect 4756 97 4828 103
rect 4932 97 5052 103
rect 5156 97 5244 103
rect 5252 97 5356 103
rect 5668 97 5724 103
rect 5764 97 5884 103
rect 6020 97 6460 103
rect 6468 97 6620 103
rect 6756 97 6924 103
rect 6948 97 7020 103
rect 7060 97 7228 103
rect 7396 97 7420 103
rect 8036 97 8076 103
rect 148 77 204 83
rect 772 77 940 83
rect 1396 77 1532 83
rect 1540 77 1564 83
rect 1572 77 1756 83
rect 1764 77 1868 83
rect 1892 77 2060 83
rect 6212 77 6316 83
rect 6324 77 7356 83
rect 1736 14 1784 16
rect 1736 6 1740 14
rect 1750 6 1756 14
rect 1764 6 1770 14
rect 1780 6 1784 14
rect 1736 4 1784 6
rect 4808 14 4856 16
rect 4808 6 4812 14
rect 4822 6 4828 14
rect 4836 6 4842 14
rect 4852 6 4856 14
rect 4808 4 4856 6
<< m4contact >>
rect 3276 5806 3278 5814
rect 3278 5806 3284 5814
rect 3292 5806 3300 5814
rect 3308 5806 3314 5814
rect 3314 5806 3316 5814
rect 6348 5806 6350 5814
rect 6350 5806 6356 5814
rect 6364 5806 6372 5814
rect 6380 5806 6386 5814
rect 6386 5806 6388 5814
rect 6204 5796 6212 5804
rect 1116 5756 1124 5764
rect 6108 5756 6116 5764
rect 860 5736 868 5744
rect 5692 5736 5700 5744
rect 7356 5736 7364 5744
rect 7644 5736 7652 5744
rect 7868 5736 7876 5744
rect 5836 5716 5844 5724
rect 8028 5716 8036 5724
rect 5692 5676 5700 5684
rect 5772 5676 5780 5684
rect 5884 5676 5892 5684
rect 1820 5656 1828 5664
rect 1564 5636 1572 5644
rect 7452 5616 7460 5624
rect 1740 5606 1742 5614
rect 1742 5606 1748 5614
rect 1756 5606 1764 5614
rect 1772 5606 1778 5614
rect 1778 5606 1780 5614
rect 4812 5606 4814 5614
rect 4814 5606 4820 5614
rect 4828 5606 4836 5614
rect 4844 5606 4850 5614
rect 4850 5606 4852 5614
rect 7420 5576 7428 5584
rect 5564 5556 5572 5564
rect 2428 5496 2436 5504
rect 2492 5496 2500 5504
rect 5884 5496 5892 5504
rect 1116 5476 1124 5484
rect 7996 5476 8004 5484
rect 8124 5476 8132 5484
rect 3836 5456 3844 5464
rect 4316 5456 4324 5464
rect 4732 5416 4740 5424
rect 3276 5406 3278 5414
rect 3278 5406 3284 5414
rect 3292 5406 3300 5414
rect 3308 5406 3314 5414
rect 3314 5406 3316 5414
rect 6348 5406 6350 5414
rect 6350 5406 6356 5414
rect 6364 5406 6372 5414
rect 6380 5406 6386 5414
rect 6386 5406 6388 5414
rect 28 5376 36 5384
rect 7772 5376 7780 5384
rect 4316 5356 4324 5364
rect 7068 5356 7076 5364
rect 5564 5336 5572 5344
rect 6108 5336 6116 5344
rect 7932 5336 7940 5344
rect 4172 5316 4180 5324
rect 4252 5316 4260 5324
rect 4732 5316 4740 5324
rect 8124 5316 8132 5324
rect 860 5296 868 5304
rect 7068 5296 7076 5304
rect 1564 5236 1572 5244
rect 4092 5236 4100 5244
rect 1740 5206 1742 5214
rect 1742 5206 1748 5214
rect 1756 5206 1764 5214
rect 1772 5206 1778 5214
rect 1778 5206 1780 5214
rect 4812 5206 4814 5214
rect 4814 5206 4820 5214
rect 4828 5206 4836 5214
rect 4844 5206 4850 5214
rect 4850 5206 4852 5214
rect 3868 5196 3876 5204
rect 3612 5136 3620 5144
rect 3228 5116 3236 5124
rect 3836 5116 3844 5124
rect 8092 5116 8100 5124
rect 3612 5096 3620 5104
rect 6908 5096 6916 5104
rect 7836 5096 7844 5104
rect 284 5076 292 5084
rect 5500 5076 5508 5084
rect 3004 5056 3012 5064
rect 7164 5056 7172 5064
rect 4188 5036 4196 5044
rect 5564 5036 5572 5044
rect 6908 5036 6916 5044
rect 7996 5036 8004 5044
rect 3868 5016 3876 5024
rect 7676 5016 7684 5024
rect 3276 5006 3278 5014
rect 3278 5006 3284 5014
rect 3292 5006 3300 5014
rect 3308 5006 3314 5014
rect 3314 5006 3316 5014
rect 6348 5006 6350 5014
rect 6350 5006 6356 5014
rect 6364 5006 6372 5014
rect 6380 5006 6386 5014
rect 6386 5006 6388 5014
rect 348 4996 356 5004
rect 4732 4996 4740 5004
rect 2876 4976 2884 4984
rect 7228 4976 7236 4984
rect 7356 4976 7364 4984
rect 7900 4976 7908 4984
rect 3004 4956 3012 4964
rect 3436 4956 3444 4964
rect 7612 4956 7620 4964
rect 284 4936 292 4944
rect 1820 4936 1828 4944
rect 7740 4936 7748 4944
rect 7996 4936 8004 4944
rect 3356 4916 3364 4924
rect 5212 4916 5220 4924
rect 7228 4916 7236 4924
rect 8124 4916 8132 4924
rect 3164 4896 3172 4904
rect 572 4876 580 4884
rect 3228 4876 3236 4884
rect 5788 4876 5796 4884
rect 3356 4856 3364 4864
rect 7644 4856 7652 4864
rect 7900 4856 7908 4864
rect 5052 4836 5060 4844
rect 4444 4816 4452 4824
rect 1740 4806 1742 4814
rect 1742 4806 1748 4814
rect 1756 4806 1764 4814
rect 1772 4806 1778 4814
rect 1778 4806 1780 4814
rect 4812 4806 4814 4814
rect 4814 4806 4820 4814
rect 4828 4806 4836 4814
rect 4844 4806 4850 4814
rect 4850 4806 4852 4814
rect 2044 4756 2052 4764
rect 7964 4756 7972 4764
rect 8060 4736 8068 4744
rect 7580 4716 7588 4724
rect 5340 4696 5348 4704
rect 5468 4696 5476 4704
rect 572 4676 580 4684
rect 7164 4656 7172 4664
rect 8060 4656 8068 4664
rect 60 4636 68 4644
rect 284 4636 292 4644
rect 2044 4636 2052 4644
rect 5340 4636 5348 4644
rect 5788 4636 5796 4644
rect 4092 4616 4100 4624
rect 4444 4616 4452 4624
rect 5052 4616 5060 4624
rect 7708 4616 7716 4624
rect 3276 4606 3278 4614
rect 3278 4606 3284 4614
rect 3292 4606 3300 4614
rect 3308 4606 3314 4614
rect 3314 4606 3316 4614
rect 6348 4606 6350 4614
rect 6350 4606 6356 4614
rect 6364 4606 6372 4614
rect 6380 4606 6386 4614
rect 6386 4606 6388 4614
rect 1468 4596 1476 4604
rect 1820 4596 1828 4604
rect 4572 4596 4580 4604
rect 348 4576 356 4584
rect 3868 4576 3876 4584
rect 7548 4596 7556 4604
rect 6492 4576 6500 4584
rect 2700 4556 2708 4564
rect 7580 4556 7588 4564
rect 2140 4536 2148 4544
rect 7612 4536 7620 4544
rect 4316 4516 4324 4524
rect 4604 4516 4612 4524
rect 7740 4516 7748 4524
rect 2140 4496 2148 4504
rect 2652 4496 2660 4504
rect 1596 4476 1604 4484
rect 7292 4476 7300 4484
rect 8124 4476 8132 4484
rect 5180 4456 5188 4464
rect 6140 4456 6148 4464
rect 2044 4436 2052 4444
rect 3164 4436 3172 4444
rect 5948 4436 5956 4444
rect 7996 4436 8004 4444
rect 3356 4416 3364 4424
rect 5052 4416 5060 4424
rect 7420 4416 7428 4424
rect 1740 4406 1742 4414
rect 1742 4406 1748 4414
rect 1756 4406 1764 4414
rect 1772 4406 1778 4414
rect 1778 4406 1780 4414
rect 4812 4406 4814 4414
rect 4814 4406 4820 4414
rect 4828 4406 4836 4414
rect 4844 4406 4850 4414
rect 4850 4406 4852 4414
rect 2428 4396 2436 4404
rect 3164 4396 3172 4404
rect 7516 4396 7524 4404
rect 2876 4376 2884 4384
rect 3868 4336 3876 4344
rect 4572 4316 4580 4324
rect 5532 4316 5540 4324
rect 7676 4316 7684 4324
rect 828 4296 836 4304
rect 3484 4296 3492 4304
rect 4988 4296 4996 4304
rect 5564 4296 5572 4304
rect 7996 4296 8004 4304
rect 8028 4296 8036 4304
rect 1436 4276 1444 4284
rect 28 4256 36 4264
rect 252 4256 260 4264
rect 860 4256 868 4264
rect 3132 4276 3140 4284
rect 5052 4276 5060 4284
rect 6300 4276 6308 4284
rect 6684 4276 6692 4284
rect 7772 4276 7780 4284
rect 4508 4256 4516 4264
rect 3164 4236 3172 4244
rect 4732 4236 4740 4244
rect 5404 4236 5412 4244
rect 7132 4236 7140 4244
rect 7708 4216 7716 4224
rect 3276 4206 3278 4214
rect 3278 4206 3284 4214
rect 3292 4206 3300 4214
rect 3308 4206 3314 4214
rect 3314 4206 3316 4214
rect 6348 4206 6350 4214
rect 6350 4206 6356 4214
rect 6364 4206 6372 4214
rect 6380 4206 6386 4214
rect 6386 4206 6388 4214
rect 188 4196 196 4204
rect 3004 4196 3012 4204
rect 4188 4196 4196 4204
rect 4508 4196 4516 4204
rect 6492 4196 6500 4204
rect 828 4176 836 4184
rect 3388 4176 3396 4184
rect 3772 4176 3780 4184
rect 5276 4176 5284 4184
rect 6140 4176 6148 4184
rect 8060 4176 8068 4184
rect 3644 4156 3652 4164
rect 5340 4156 5348 4164
rect 7900 4156 7908 4164
rect 8124 4156 8132 4164
rect 3772 4136 3780 4144
rect 4892 4136 4900 4144
rect 6684 4136 6692 4144
rect 7516 4136 7524 4144
rect 1436 4116 1444 4124
rect 2828 4116 2836 4124
rect 3676 4116 3684 4124
rect 4540 4116 4548 4124
rect 4988 4116 4996 4124
rect 2780 4096 2788 4104
rect 5276 4116 5284 4124
rect 6300 4116 6308 4124
rect 2844 4076 2852 4084
rect 3484 4076 3492 4084
rect 7804 4076 7812 4084
rect 2492 4056 2500 4064
rect 2684 4056 2692 4064
rect 5180 4056 5188 4064
rect 7740 4056 7748 4064
rect 3676 4036 3684 4044
rect 5916 4036 5924 4044
rect 6204 4036 6212 4044
rect 2844 4016 2852 4024
rect 5052 4016 5060 4024
rect 1740 4006 1742 4014
rect 1742 4006 1748 4014
rect 1756 4006 1764 4014
rect 1772 4006 1778 4014
rect 1778 4006 1780 4014
rect 4812 4006 4814 4014
rect 4814 4006 4820 4014
rect 4828 4006 4836 4014
rect 4844 4006 4850 4014
rect 4850 4006 4852 4014
rect 2716 3996 2724 4004
rect 3772 3996 3780 4004
rect 5500 3996 5508 4004
rect 6108 3996 6116 4004
rect 860 3976 868 3984
rect 3484 3976 3492 3984
rect 6908 3936 6916 3944
rect 7452 3936 7460 3944
rect 7676 3936 7684 3944
rect 1884 3916 1892 3924
rect 3612 3916 3620 3924
rect 3484 3876 3492 3884
rect 3548 3876 3556 3884
rect 3708 3876 3716 3884
rect 5948 3896 5956 3904
rect 6620 3896 6628 3904
rect 7964 3896 7972 3904
rect 6236 3876 6244 3884
rect 7292 3876 7300 3884
rect 3612 3856 3620 3864
rect 3740 3856 3748 3864
rect 7900 3856 7908 3864
rect 1468 3816 1476 3824
rect 3548 3816 3556 3824
rect 4540 3816 4548 3824
rect 4892 3816 4900 3824
rect 3276 3806 3278 3814
rect 3278 3806 3284 3814
rect 3292 3806 3300 3814
rect 3308 3806 3314 3814
rect 3314 3806 3316 3814
rect 6348 3806 6350 3814
rect 6350 3806 6356 3814
rect 6364 3806 6372 3814
rect 6380 3806 6386 3814
rect 6386 3806 6388 3814
rect 188 3776 196 3784
rect 3740 3776 3748 3784
rect 4412 3776 4420 3784
rect 5468 3776 5476 3784
rect 6620 3796 6628 3804
rect 6428 3776 6436 3784
rect 8124 3776 8132 3784
rect 1884 3756 1892 3764
rect 4572 3756 4580 3764
rect 5500 3756 5508 3764
rect 5532 3756 5540 3764
rect 6492 3756 6500 3764
rect 7036 3756 7044 3764
rect 7804 3756 7812 3764
rect 1084 3716 1092 3724
rect 6620 3716 6628 3724
rect 7964 3716 7972 3724
rect 4572 3696 4580 3704
rect 7132 3696 7140 3704
rect 3708 3676 3716 3684
rect 6268 3676 6276 3684
rect 3932 3656 3940 3664
rect 4924 3656 4932 3664
rect 4700 3636 4708 3644
rect 4732 3636 4740 3644
rect 4988 3636 4996 3644
rect 6620 3636 6628 3644
rect 5884 3616 5892 3624
rect 1740 3606 1742 3614
rect 1742 3606 1748 3614
rect 1756 3606 1764 3614
rect 1772 3606 1778 3614
rect 1778 3606 1780 3614
rect 4812 3606 4814 3614
rect 4814 3606 4820 3614
rect 4828 3606 4836 3614
rect 4844 3606 4850 3614
rect 4850 3606 4852 3614
rect 4636 3596 4644 3604
rect 5340 3596 5348 3604
rect 5372 3596 5380 3604
rect 6140 3576 6148 3584
rect 3964 3556 3972 3564
rect 4540 3536 4548 3544
rect 5404 3536 5412 3544
rect 6972 3556 6980 3564
rect 8092 3556 8100 3564
rect 508 3516 516 3524
rect 1244 3516 1252 3524
rect 2716 3496 2724 3504
rect 5148 3496 5156 3504
rect 6492 3496 6500 3504
rect 3356 3476 3364 3484
rect 4540 3476 4548 3484
rect 7388 3476 7396 3484
rect 316 3456 324 3464
rect 6076 3456 6084 3464
rect 540 3436 548 3444
rect 2012 3436 2020 3444
rect 3676 3436 3684 3444
rect 7548 3436 7556 3444
rect 1244 3416 1252 3424
rect 1980 3416 1988 3424
rect 6108 3416 6116 3424
rect 3276 3406 3278 3414
rect 3278 3406 3284 3414
rect 3292 3406 3300 3414
rect 3308 3406 3314 3414
rect 3314 3406 3316 3414
rect 6348 3406 6350 3414
rect 6350 3406 6356 3414
rect 6364 3406 6372 3414
rect 6380 3406 6386 3414
rect 6386 3406 6388 3414
rect 508 3396 516 3404
rect 3356 3396 3364 3404
rect 5148 3396 5156 3404
rect 412 3376 420 3384
rect 3612 3376 3620 3384
rect 5468 3376 5476 3384
rect 7772 3376 7780 3384
rect 732 3356 740 3364
rect 252 3336 260 3344
rect 1532 3336 1540 3344
rect 3100 3336 3108 3344
rect 3676 3336 3684 3344
rect 4636 3336 4644 3344
rect 6076 3336 6084 3344
rect 6908 3336 6916 3344
rect 7452 3336 7460 3344
rect 4284 3316 4292 3324
rect 5084 3316 5092 3324
rect 5212 3296 5220 3304
rect 7708 3296 7716 3304
rect 8028 3296 8036 3304
rect 3612 3276 3620 3284
rect 5084 3276 5092 3284
rect 1532 3256 1540 3264
rect 1980 3236 1988 3244
rect 2812 3236 2820 3244
rect 7292 3236 7300 3244
rect 1740 3206 1742 3214
rect 1742 3206 1748 3214
rect 1756 3206 1764 3214
rect 1772 3206 1778 3214
rect 1778 3206 1780 3214
rect 4812 3206 4814 3214
rect 4814 3206 4820 3214
rect 4828 3206 4836 3214
rect 4844 3206 4850 3214
rect 4850 3206 4852 3214
rect 3772 3196 3780 3204
rect 540 3176 548 3184
rect 4060 3176 4068 3184
rect 4892 3176 4900 3184
rect 6236 3176 6244 3184
rect 6460 3176 6468 3184
rect 7516 3176 7524 3184
rect 1084 3156 1092 3164
rect 2460 3136 2468 3144
rect 3644 3116 3652 3124
rect 6652 3116 6660 3124
rect 316 3096 324 3104
rect 7772 3096 7780 3104
rect 7868 3096 7876 3104
rect 1372 3076 1380 3084
rect 4412 3076 4420 3084
rect 6268 3076 6276 3084
rect 7292 3076 7300 3084
rect 3036 3056 3044 3064
rect 4668 3056 4676 3064
rect 6652 3056 6660 3064
rect 60 3036 68 3044
rect 4060 3036 4068 3044
rect 4540 3036 4548 3044
rect 7708 3016 7716 3024
rect 7772 3016 7780 3024
rect 3276 3006 3278 3014
rect 3278 3006 3284 3014
rect 3292 3006 3300 3014
rect 3308 3006 3314 3014
rect 3314 3006 3316 3014
rect 6348 3006 6350 3014
rect 6350 3006 6356 3014
rect 6364 3006 6372 3014
rect 6380 3006 6386 3014
rect 6386 3006 6388 3014
rect 6428 2996 6436 3004
rect 5564 2976 5572 2984
rect 988 2956 996 2964
rect 3644 2956 3652 2964
rect 7388 2956 7396 2964
rect 2460 2916 2468 2924
rect 3196 2916 3204 2924
rect 3388 2916 3396 2924
rect 3644 2916 3652 2924
rect 5148 2916 5156 2924
rect 8028 2916 8036 2924
rect 4892 2896 4900 2904
rect 7292 2896 7300 2904
rect 7996 2876 8004 2884
rect 2108 2856 2116 2864
rect 3164 2856 3172 2864
rect 7836 2856 7844 2864
rect 1532 2836 1540 2844
rect 2812 2836 2820 2844
rect 3676 2836 3684 2844
rect 5052 2836 5060 2844
rect 5436 2836 5444 2844
rect 6140 2816 6148 2824
rect 1740 2806 1742 2814
rect 1742 2806 1748 2814
rect 1756 2806 1764 2814
rect 1772 2806 1778 2814
rect 1778 2806 1780 2814
rect 4812 2806 4814 2814
rect 4814 2806 4820 2814
rect 4828 2806 4836 2814
rect 4844 2806 4850 2814
rect 4850 2806 4852 2814
rect 3132 2796 3140 2804
rect 4636 2796 4644 2804
rect 4700 2796 4708 2804
rect 5884 2796 5892 2804
rect 7068 2796 7076 2804
rect 8028 2776 8036 2784
rect 412 2756 420 2764
rect 6300 2736 6308 2744
rect 5948 2716 5956 2724
rect 7932 2716 7940 2724
rect 860 2676 868 2684
rect 2524 2696 2532 2704
rect 2684 2696 2692 2704
rect 2140 2676 2148 2684
rect 3100 2676 3108 2684
rect 4668 2676 4676 2684
rect 6684 2676 6692 2684
rect 8060 2676 8068 2684
rect 4540 2656 4548 2664
rect 6268 2656 6276 2664
rect 5148 2636 5156 2644
rect 6204 2616 6212 2624
rect 6236 2616 6244 2624
rect 3276 2606 3278 2614
rect 3278 2606 3284 2614
rect 3292 2606 3300 2614
rect 3308 2606 3314 2614
rect 3314 2606 3316 2614
rect 6348 2606 6350 2614
rect 6350 2606 6356 2614
rect 6364 2606 6372 2614
rect 6380 2606 6386 2614
rect 6386 2606 6388 2614
rect 3100 2596 3108 2604
rect 4220 2596 4228 2604
rect 4252 2596 4260 2604
rect 8060 2596 8068 2604
rect 4188 2556 4196 2564
rect 4220 2556 4228 2564
rect 4604 2536 4612 2544
rect 6268 2516 6276 2524
rect 6428 2516 6436 2524
rect 6620 2516 6628 2524
rect 3644 2496 3652 2504
rect 5564 2496 5572 2504
rect 7740 2496 7748 2504
rect 7804 2496 7812 2504
rect 4700 2476 4708 2484
rect 5372 2476 5380 2484
rect 4284 2456 4292 2464
rect 4988 2436 4996 2444
rect 7580 2436 7588 2444
rect 4316 2416 4324 2424
rect 4412 2416 4420 2424
rect 1740 2406 1742 2414
rect 1742 2406 1748 2414
rect 1756 2406 1764 2414
rect 1772 2406 1778 2414
rect 1778 2406 1780 2414
rect 4812 2406 4814 2414
rect 4814 2406 4820 2414
rect 4828 2406 4836 2414
rect 4844 2406 4850 2414
rect 4850 2406 4852 2414
rect 5948 2396 5956 2404
rect 3164 2376 3172 2384
rect 3356 2376 3364 2384
rect 4060 2376 4068 2384
rect 3996 2356 4004 2364
rect 4764 2356 4772 2364
rect 5916 2356 5924 2364
rect 6844 2356 6852 2364
rect 7036 2356 7044 2364
rect 6140 2336 6148 2344
rect 6460 2336 6468 2344
rect 3068 2316 3076 2324
rect 3964 2316 3972 2324
rect 4764 2316 4772 2324
rect 2012 2296 2020 2304
rect 2780 2296 2788 2304
rect 4252 2296 4260 2304
rect 1596 2276 1604 2284
rect 2428 2276 2436 2284
rect 2748 2276 2756 2284
rect 3036 2276 3044 2284
rect 4188 2276 4196 2284
rect 7676 2276 7684 2284
rect 2556 2256 2564 2264
rect 2716 2256 2724 2264
rect 3388 2256 3396 2264
rect 5692 2236 5700 2244
rect 6716 2236 6724 2244
rect 7356 2216 7364 2224
rect 3276 2206 3278 2214
rect 3278 2206 3284 2214
rect 3292 2206 3300 2214
rect 3308 2206 3314 2214
rect 3314 2206 3316 2214
rect 6348 2206 6350 2214
rect 6350 2206 6356 2214
rect 6364 2206 6372 2214
rect 6380 2206 6386 2214
rect 6386 2206 6388 2214
rect 2780 2176 2788 2184
rect 3932 2196 3940 2204
rect 4700 2176 4708 2184
rect 7580 2176 7588 2184
rect 732 2156 740 2164
rect 2108 2156 2116 2164
rect 2716 2156 2724 2164
rect 4668 2156 4676 2164
rect 6300 2156 6308 2164
rect 988 2136 996 2144
rect 4188 2136 4196 2144
rect 4316 2136 4324 2144
rect 6204 2136 6212 2144
rect 6236 2136 6244 2144
rect 1820 2116 1828 2124
rect 2748 2116 2756 2124
rect 2780 2096 2788 2104
rect 7708 2096 7716 2104
rect 7772 2096 7780 2104
rect 3996 2056 4004 2064
rect 4540 2016 4548 2024
rect 4636 2016 4644 2024
rect 1740 2006 1742 2014
rect 1742 2006 1748 2014
rect 1756 2006 1764 2014
rect 1772 2006 1778 2014
rect 1778 2006 1780 2014
rect 4812 2006 4814 2014
rect 4814 2006 4820 2014
rect 4828 2006 4836 2014
rect 4844 2006 4850 2014
rect 4850 2006 4852 2014
rect 1372 1996 1380 2004
rect 3100 1996 3108 2004
rect 3196 1996 3204 2004
rect 5436 1976 5444 1984
rect 220 1956 228 1964
rect 2844 1956 2852 1964
rect 3388 1956 3396 1964
rect 7452 1956 7460 1964
rect 220 1916 228 1924
rect 1372 1916 1380 1924
rect 6844 1916 6852 1924
rect 4412 1896 4420 1904
rect 4604 1896 4612 1904
rect 5564 1896 5572 1904
rect 5692 1896 5700 1904
rect 7452 1896 7460 1904
rect 3964 1876 3972 1884
rect 2876 1836 2884 1844
rect 2780 1816 2788 1824
rect 3356 1816 3364 1824
rect 3276 1806 3278 1814
rect 3278 1806 3284 1814
rect 3292 1806 3300 1814
rect 3308 1806 3314 1814
rect 3314 1806 3316 1814
rect 4604 1796 4612 1804
rect 5692 1816 5700 1824
rect 6348 1806 6350 1814
rect 6350 1806 6356 1814
rect 6364 1806 6372 1814
rect 6380 1806 6386 1814
rect 6386 1806 6388 1814
rect 1180 1776 1188 1784
rect 2108 1776 2116 1784
rect 3772 1776 3780 1784
rect 2876 1756 2884 1764
rect 6140 1776 6148 1784
rect 6524 1776 6532 1784
rect 4476 1756 4484 1764
rect 7516 1756 7524 1764
rect 2044 1736 2052 1744
rect 2844 1736 2852 1744
rect 3420 1736 3428 1744
rect 4412 1736 4420 1744
rect 6236 1736 6244 1744
rect 4092 1716 4100 1724
rect 5692 1716 5700 1724
rect 3772 1696 3780 1704
rect 3420 1676 3428 1684
rect 4508 1696 4516 1704
rect 4380 1656 4388 1664
rect 4412 1656 4420 1664
rect 2524 1636 2532 1644
rect 700 1616 708 1624
rect 4508 1616 4516 1624
rect 1740 1606 1742 1614
rect 1742 1606 1748 1614
rect 1756 1606 1764 1614
rect 1772 1606 1778 1614
rect 1778 1606 1780 1614
rect 4812 1606 4814 1614
rect 4814 1606 4820 1614
rect 4828 1606 4836 1614
rect 4844 1606 4850 1614
rect 4850 1606 4852 1614
rect 3004 1576 3012 1584
rect 5084 1576 5092 1584
rect 6524 1536 6532 1544
rect 2300 1516 2308 1524
rect 3068 1496 3076 1504
rect 3452 1496 3460 1504
rect 5820 1496 5828 1504
rect 6428 1496 6436 1504
rect 6716 1516 6724 1524
rect 6972 1496 6980 1504
rect 700 1476 708 1484
rect 7420 1476 7428 1484
rect 6748 1456 6756 1464
rect 7356 1456 7364 1464
rect 4092 1416 4100 1424
rect 4540 1416 4548 1424
rect 5948 1416 5956 1424
rect 6972 1416 6980 1424
rect 3276 1406 3278 1414
rect 3278 1406 3284 1414
rect 3292 1406 3300 1414
rect 3308 1406 3314 1414
rect 3314 1406 3316 1414
rect 6348 1406 6350 1414
rect 6350 1406 6356 1414
rect 6364 1406 6372 1414
rect 6380 1406 6386 1414
rect 6386 1406 6388 1414
rect 7068 1396 7076 1404
rect 2428 1356 2436 1364
rect 5916 1356 5924 1364
rect 6236 1336 6244 1344
rect 2652 1296 2660 1304
rect 5820 1296 5828 1304
rect 4924 1276 4932 1284
rect 1740 1206 1742 1214
rect 1742 1206 1748 1214
rect 1756 1206 1764 1214
rect 1772 1206 1778 1214
rect 1778 1206 1780 1214
rect 4812 1206 4814 1214
rect 4814 1206 4820 1214
rect 4828 1206 4836 1214
rect 4844 1206 4850 1214
rect 4850 1206 4852 1214
rect 3356 1196 3364 1204
rect 604 1176 612 1184
rect 4252 1176 4260 1184
rect 5948 1176 5956 1184
rect 412 1096 420 1104
rect 1372 1096 1380 1104
rect 2108 1096 2116 1104
rect 3708 1096 3716 1104
rect 3868 1096 3876 1104
rect 5084 1096 5092 1104
rect 636 1076 644 1084
rect 1180 1076 1188 1084
rect 2684 1076 2692 1084
rect 6748 1076 6756 1084
rect 2044 1056 2052 1064
rect 3676 1056 3684 1064
rect 3932 1056 3940 1064
rect 4348 1056 4356 1064
rect 1404 1016 1412 1024
rect 2556 1016 2564 1024
rect 3100 1016 3108 1024
rect 3932 1016 3940 1024
rect 3276 1006 3278 1014
rect 3278 1006 3284 1014
rect 3292 1006 3300 1014
rect 3308 1006 3314 1014
rect 3314 1006 3316 1014
rect 6348 1006 6350 1014
rect 6350 1006 6356 1014
rect 6364 1006 6372 1014
rect 6380 1006 6386 1014
rect 6386 1006 6388 1014
rect 1436 996 1444 1004
rect 1532 996 1540 1004
rect 3004 996 3012 1004
rect 4348 996 4356 1004
rect 5468 976 5476 984
rect 5916 976 5924 984
rect 348 936 356 944
rect 3676 936 3684 944
rect 5084 936 5092 944
rect 6108 936 6116 944
rect 1212 916 1220 924
rect 1404 916 1412 924
rect 1436 916 1444 924
rect 4348 916 4356 924
rect 1596 896 1604 904
rect 1372 856 1380 864
rect 7612 836 7620 844
rect 7708 836 7716 844
rect 2684 816 2692 824
rect 5564 816 5572 824
rect 1740 806 1742 814
rect 1742 806 1748 814
rect 1756 806 1764 814
rect 1772 806 1778 814
rect 1778 806 1780 814
rect 4812 806 4814 814
rect 4814 806 4820 814
rect 4828 806 4836 814
rect 4844 806 4850 814
rect 4850 806 4852 814
rect 604 776 612 784
rect 4476 776 4484 784
rect 4252 756 4260 764
rect 3708 736 3716 744
rect 8060 736 8068 744
rect 3868 716 3876 724
rect 1532 696 1540 704
rect 3708 696 3716 704
rect 7900 696 7908 704
rect 4380 676 4388 684
rect 4700 676 4708 684
rect 7804 676 7812 684
rect 3452 656 3460 664
rect 3964 656 3972 664
rect 6076 656 6084 664
rect 1212 616 1220 624
rect 1596 616 1604 624
rect 4700 616 4708 624
rect 3276 606 3278 614
rect 3278 606 3284 614
rect 3292 606 3300 614
rect 3308 606 3314 614
rect 3314 606 3316 614
rect 6348 606 6350 614
rect 6350 606 6356 614
rect 6364 606 6372 614
rect 6380 606 6386 614
rect 6386 606 6388 614
rect 1212 576 1220 584
rect 2652 576 2660 584
rect 636 556 644 564
rect 188 536 196 544
rect 6076 516 6084 524
rect 8060 516 8068 524
rect 348 496 356 504
rect 3580 476 3588 484
rect 8028 476 8036 484
rect 412 456 420 464
rect 2300 456 2308 464
rect 3356 436 3364 444
rect 4476 436 4484 444
rect 1740 406 1742 414
rect 1742 406 1748 414
rect 1756 406 1764 414
rect 1772 406 1778 414
rect 1778 406 1780 414
rect 4812 406 4814 414
rect 4814 406 4820 414
rect 4828 406 4836 414
rect 4844 406 4850 414
rect 4850 406 4852 414
rect 3228 376 3236 384
rect 2716 316 2724 324
rect 7900 316 7908 324
rect 7964 316 7972 324
rect 5468 296 5476 304
rect 2716 276 2724 284
rect 3740 276 3748 284
rect 6108 276 6116 284
rect 7420 276 7428 284
rect 7964 256 7972 264
rect 3580 236 3588 244
rect 7612 236 7620 244
rect 8060 236 8068 244
rect 188 216 196 224
rect 3276 206 3278 214
rect 3278 206 3284 214
rect 3292 206 3300 214
rect 3308 206 3314 214
rect 3314 206 3316 214
rect 6348 206 6350 214
rect 6350 206 6356 214
rect 6364 206 6372 214
rect 6380 206 6386 214
rect 6386 206 6388 214
rect 5724 196 5732 204
rect 2076 176 2084 184
rect 3740 176 3748 184
rect 2140 156 2148 164
rect 3228 136 3236 144
rect 5564 156 5572 164
rect 5724 136 5732 144
rect 6556 136 6564 144
rect 6652 136 6660 144
rect 7868 156 7876 164
rect 6876 116 6884 124
rect 7868 116 7876 124
rect 6940 96 6948 104
rect 1740 6 1742 14
rect 1742 6 1748 14
rect 1756 6 1764 14
rect 1772 6 1778 14
rect 1778 6 1780 14
rect 4812 6 4814 14
rect 4814 6 4820 14
rect 4828 6 4836 14
rect 4844 6 4850 14
rect 4850 6 4852 14
<< metal4 >>
rect 1114 5764 1126 5766
rect 1114 5756 1116 5764
rect 1124 5756 1126 5764
rect 858 5744 870 5746
rect 858 5736 860 5744
rect 868 5736 870 5744
rect 26 5384 38 5386
rect 26 5376 28 5384
rect 36 5376 38 5384
rect 26 4264 38 5376
rect 858 5304 870 5736
rect 1114 5484 1126 5756
rect 1114 5476 1116 5484
rect 1124 5476 1126 5484
rect 1114 5474 1126 5476
rect 1562 5644 1574 5646
rect 1562 5636 1564 5644
rect 1572 5636 1574 5644
rect 858 5296 860 5304
rect 868 5296 870 5304
rect 858 5294 870 5296
rect 1562 5244 1574 5636
rect 1562 5236 1564 5244
rect 1572 5236 1574 5244
rect 1562 5234 1574 5236
rect 1736 5614 1784 5840
rect 3272 5814 3320 5840
rect 3272 5806 3276 5814
rect 3284 5806 3292 5814
rect 3300 5806 3308 5814
rect 3316 5806 3320 5814
rect 1736 5606 1740 5614
rect 1748 5606 1756 5614
rect 1764 5606 1772 5614
rect 1780 5606 1784 5614
rect 1736 5214 1784 5606
rect 1736 5206 1740 5214
rect 1748 5206 1756 5214
rect 1764 5206 1772 5214
rect 1780 5206 1784 5214
rect 282 5084 294 5086
rect 282 5076 284 5084
rect 292 5076 294 5084
rect 282 4944 294 5076
rect 282 4936 284 4944
rect 292 4936 294 4944
rect 26 4256 28 4264
rect 36 4256 38 4264
rect 26 4254 38 4256
rect 58 4644 70 4646
rect 58 4636 60 4644
rect 68 4636 70 4644
rect 58 3044 70 4636
rect 282 4644 294 4936
rect 282 4636 284 4644
rect 292 4636 294 4644
rect 282 4634 294 4636
rect 346 5004 358 5006
rect 346 4996 348 5004
rect 356 4996 358 5004
rect 346 4584 358 4996
rect 570 4884 582 4886
rect 570 4876 572 4884
rect 580 4876 582 4884
rect 570 4684 582 4876
rect 570 4676 572 4684
rect 580 4676 582 4684
rect 570 4674 582 4676
rect 1736 4814 1784 5206
rect 1818 5664 1830 5666
rect 1818 5656 1820 5664
rect 1828 5656 1830 5664
rect 1818 4944 1830 5656
rect 1818 4936 1820 4944
rect 1828 4936 1830 4944
rect 1818 4934 1830 4936
rect 2426 5504 2438 5506
rect 2426 5496 2428 5504
rect 2436 5496 2438 5504
rect 1736 4806 1740 4814
rect 1748 4806 1756 4814
rect 1764 4806 1772 4814
rect 1780 4806 1784 4814
rect 346 4576 348 4584
rect 356 4576 358 4584
rect 346 4574 358 4576
rect 1466 4604 1478 4606
rect 1466 4596 1468 4604
rect 1476 4596 1478 4604
rect 826 4304 838 4306
rect 826 4296 828 4304
rect 836 4296 838 4304
rect 250 4264 262 4266
rect 250 4256 252 4264
rect 260 4256 262 4264
rect 186 4204 198 4206
rect 186 4196 188 4204
rect 196 4196 198 4204
rect 186 3784 198 4196
rect 186 3776 188 3784
rect 196 3776 198 3784
rect 186 3774 198 3776
rect 250 3344 262 4256
rect 826 4184 838 4296
rect 1434 4284 1446 4286
rect 1434 4276 1436 4284
rect 1444 4276 1446 4284
rect 826 4176 828 4184
rect 836 4176 838 4184
rect 826 4174 838 4176
rect 858 4264 870 4266
rect 858 4256 860 4264
rect 868 4256 870 4264
rect 858 3984 870 4256
rect 1434 4124 1446 4276
rect 1434 4116 1436 4124
rect 1444 4116 1446 4124
rect 1434 4114 1446 4116
rect 858 3976 860 3984
rect 868 3976 870 3984
rect 506 3524 518 3526
rect 506 3516 508 3524
rect 516 3516 518 3524
rect 250 3336 252 3344
rect 260 3336 262 3344
rect 250 3334 262 3336
rect 314 3464 326 3466
rect 314 3456 316 3464
rect 324 3456 326 3464
rect 314 3104 326 3456
rect 506 3404 518 3516
rect 506 3396 508 3404
rect 516 3396 518 3404
rect 506 3394 518 3396
rect 538 3444 550 3446
rect 538 3436 540 3444
rect 548 3436 550 3444
rect 314 3096 316 3104
rect 324 3096 326 3104
rect 314 3094 326 3096
rect 410 3384 422 3386
rect 410 3376 412 3384
rect 420 3376 422 3384
rect 58 3036 60 3044
rect 68 3036 70 3044
rect 58 3034 70 3036
rect 410 2764 422 3376
rect 538 3184 550 3436
rect 538 3176 540 3184
rect 548 3176 550 3184
rect 538 3174 550 3176
rect 730 3364 742 3366
rect 730 3356 732 3364
rect 740 3356 742 3364
rect 410 2756 412 2764
rect 420 2756 422 2764
rect 410 2754 422 2756
rect 730 2164 742 3356
rect 858 2684 870 3976
rect 1466 3824 1478 4596
rect 1466 3816 1468 3824
rect 1476 3816 1478 3824
rect 1466 3814 1478 3816
rect 1594 4484 1606 4486
rect 1594 4476 1596 4484
rect 1604 4476 1606 4484
rect 1082 3724 1094 3726
rect 1082 3716 1084 3724
rect 1092 3716 1094 3724
rect 1082 3164 1094 3716
rect 1242 3524 1254 3526
rect 1242 3516 1244 3524
rect 1252 3516 1254 3524
rect 1242 3424 1254 3516
rect 1242 3416 1244 3424
rect 1252 3416 1254 3424
rect 1242 3414 1254 3416
rect 1082 3156 1084 3164
rect 1092 3156 1094 3164
rect 1082 3154 1094 3156
rect 1530 3344 1542 3346
rect 1530 3336 1532 3344
rect 1540 3336 1542 3344
rect 1530 3264 1542 3336
rect 1530 3256 1532 3264
rect 1540 3256 1542 3264
rect 1370 3084 1382 3086
rect 1370 3076 1372 3084
rect 1380 3076 1382 3084
rect 858 2676 860 2684
rect 868 2676 870 2684
rect 858 2674 870 2676
rect 986 2964 998 2966
rect 986 2956 988 2964
rect 996 2956 998 2964
rect 730 2156 732 2164
rect 740 2156 742 2164
rect 730 2154 742 2156
rect 986 2144 998 2956
rect 986 2136 988 2144
rect 996 2136 998 2144
rect 986 2134 998 2136
rect 1370 2004 1382 3076
rect 1530 2844 1542 3256
rect 1530 2836 1532 2844
rect 1540 2836 1542 2844
rect 1530 2834 1542 2836
rect 1594 2284 1606 4476
rect 1594 2276 1596 2284
rect 1604 2276 1606 2284
rect 1594 2274 1606 2276
rect 1736 4414 1784 4806
rect 2042 4764 2054 4766
rect 2042 4756 2044 4764
rect 2052 4756 2054 4764
rect 2042 4644 2054 4756
rect 2042 4636 2044 4644
rect 2052 4636 2054 4644
rect 1736 4406 1740 4414
rect 1748 4406 1756 4414
rect 1764 4406 1772 4414
rect 1780 4406 1784 4414
rect 1736 4014 1784 4406
rect 1736 4006 1740 4014
rect 1748 4006 1756 4014
rect 1764 4006 1772 4014
rect 1780 4006 1784 4014
rect 1736 3614 1784 4006
rect 1736 3606 1740 3614
rect 1748 3606 1756 3614
rect 1764 3606 1772 3614
rect 1780 3606 1784 3614
rect 1736 3214 1784 3606
rect 1736 3206 1740 3214
rect 1748 3206 1756 3214
rect 1764 3206 1772 3214
rect 1780 3206 1784 3214
rect 1736 2814 1784 3206
rect 1736 2806 1740 2814
rect 1748 2806 1756 2814
rect 1764 2806 1772 2814
rect 1780 2806 1784 2814
rect 1736 2414 1784 2806
rect 1736 2406 1740 2414
rect 1748 2406 1756 2414
rect 1764 2406 1772 2414
rect 1780 2406 1784 2414
rect 1370 1996 1372 2004
rect 1380 1996 1382 2004
rect 1370 1994 1382 1996
rect 1736 2014 1784 2406
rect 1818 4604 1830 4606
rect 1818 4596 1820 4604
rect 1828 4596 1830 4604
rect 1818 2124 1830 4596
rect 2042 4444 2054 4636
rect 2042 4436 2044 4444
rect 2052 4436 2054 4444
rect 2042 4434 2054 4436
rect 2138 4544 2150 4546
rect 2138 4536 2140 4544
rect 2148 4536 2150 4544
rect 2138 4504 2150 4536
rect 2138 4496 2140 4504
rect 2148 4496 2150 4504
rect 1882 3924 1894 3926
rect 1882 3916 1884 3924
rect 1892 3916 1894 3924
rect 1882 3764 1894 3916
rect 1882 3756 1884 3764
rect 1892 3756 1894 3764
rect 1882 3754 1894 3756
rect 2010 3444 2022 3446
rect 2010 3436 2012 3444
rect 2020 3436 2022 3444
rect 1978 3424 1990 3426
rect 1978 3416 1980 3424
rect 1988 3416 1990 3424
rect 1978 3244 1990 3416
rect 1978 3236 1980 3244
rect 1988 3236 1990 3244
rect 1978 3234 1990 3236
rect 2010 2304 2022 3436
rect 2010 2296 2012 2304
rect 2020 2296 2022 2304
rect 2010 2294 2022 2296
rect 2106 2864 2118 2866
rect 2106 2856 2108 2864
rect 2116 2856 2118 2864
rect 2106 2164 2118 2856
rect 2138 2684 2150 4496
rect 2426 4404 2438 5496
rect 2426 4396 2428 4404
rect 2436 4396 2438 4404
rect 2426 4394 2438 4396
rect 2490 5504 2502 5506
rect 2490 5496 2492 5504
rect 2500 5496 2502 5504
rect 2490 4064 2502 5496
rect 3272 5414 3320 5806
rect 4808 5614 4856 5840
rect 6344 5814 6392 5840
rect 6344 5806 6348 5814
rect 6356 5806 6364 5814
rect 6372 5806 6380 5814
rect 6388 5806 6392 5814
rect 6202 5804 6214 5806
rect 6202 5796 6204 5804
rect 6212 5796 6214 5804
rect 6106 5764 6118 5766
rect 6106 5756 6108 5764
rect 6116 5756 6118 5764
rect 5690 5744 5702 5746
rect 5690 5736 5692 5744
rect 5700 5736 5702 5744
rect 5690 5684 5702 5736
rect 5818 5724 5846 5726
rect 5818 5716 5836 5724
rect 5844 5716 5846 5724
rect 5818 5714 5846 5716
rect 5818 5686 5830 5714
rect 5690 5676 5692 5684
rect 5700 5676 5702 5684
rect 5690 5674 5702 5676
rect 5770 5684 5830 5686
rect 5770 5676 5772 5684
rect 5780 5676 5830 5684
rect 5770 5674 5830 5676
rect 5882 5684 5894 5686
rect 5882 5676 5884 5684
rect 5892 5676 5894 5684
rect 4808 5606 4812 5614
rect 4820 5606 4828 5614
rect 4836 5606 4844 5614
rect 4852 5606 4856 5614
rect 3272 5406 3276 5414
rect 3284 5406 3292 5414
rect 3300 5406 3308 5414
rect 3316 5406 3320 5414
rect 3226 5124 3238 5126
rect 3226 5116 3228 5124
rect 3236 5116 3238 5124
rect 3002 5064 3014 5066
rect 3002 5056 3004 5064
rect 3012 5056 3014 5064
rect 2874 4984 2886 4986
rect 2874 4976 2876 4984
rect 2884 4976 2886 4984
rect 2650 4564 2710 4566
rect 2650 4556 2700 4564
rect 2708 4556 2710 4564
rect 2650 4554 2710 4556
rect 2650 4504 2662 4554
rect 2650 4496 2652 4504
rect 2660 4496 2662 4504
rect 2650 4494 2662 4496
rect 2874 4384 2886 4976
rect 2874 4376 2876 4384
rect 2884 4376 2886 4384
rect 2874 4374 2886 4376
rect 3002 4964 3014 5056
rect 3002 4956 3004 4964
rect 3012 4956 3014 4964
rect 3002 4204 3014 4956
rect 3162 4904 3174 4906
rect 3162 4896 3164 4904
rect 3172 4896 3174 4904
rect 3162 4444 3174 4896
rect 3226 4884 3238 5116
rect 3226 4876 3228 4884
rect 3236 4876 3238 4884
rect 3226 4874 3238 4876
rect 3272 5014 3320 5406
rect 3834 5464 3846 5466
rect 3834 5456 3836 5464
rect 3844 5456 3846 5464
rect 3610 5144 3622 5146
rect 3610 5136 3612 5144
rect 3620 5136 3622 5144
rect 3610 5104 3622 5136
rect 3834 5124 3846 5456
rect 4314 5464 4326 5466
rect 4314 5456 4316 5464
rect 4324 5456 4326 5464
rect 4314 5364 4326 5456
rect 4314 5356 4316 5364
rect 4324 5356 4326 5364
rect 4170 5324 4262 5326
rect 4170 5316 4172 5324
rect 4180 5316 4252 5324
rect 4260 5316 4262 5324
rect 4170 5314 4262 5316
rect 4090 5244 4102 5246
rect 4090 5236 4092 5244
rect 4100 5236 4102 5244
rect 3834 5116 3836 5124
rect 3844 5116 3846 5124
rect 3834 5114 3846 5116
rect 3866 5204 3878 5206
rect 3866 5196 3868 5204
rect 3876 5196 3878 5204
rect 3610 5096 3612 5104
rect 3620 5096 3622 5104
rect 3610 5094 3622 5096
rect 3866 5024 3878 5196
rect 3866 5016 3868 5024
rect 3876 5016 3878 5024
rect 3866 5014 3878 5016
rect 3272 5006 3276 5014
rect 3284 5006 3292 5014
rect 3300 5006 3308 5014
rect 3316 5006 3320 5014
rect 3162 4436 3164 4444
rect 3172 4436 3174 4444
rect 3162 4434 3174 4436
rect 3272 4614 3320 5006
rect 3354 4964 3446 4966
rect 3354 4956 3436 4964
rect 3444 4956 3446 4964
rect 3354 4954 3446 4956
rect 3354 4924 3366 4954
rect 3354 4916 3356 4924
rect 3364 4916 3366 4924
rect 3354 4914 3366 4916
rect 3272 4606 3276 4614
rect 3284 4606 3292 4614
rect 3300 4606 3308 4614
rect 3316 4606 3320 4614
rect 3162 4404 3174 4406
rect 3162 4396 3164 4404
rect 3172 4396 3174 4404
rect 3002 4196 3004 4204
rect 3012 4196 3014 4204
rect 3002 4194 3014 4196
rect 3130 4284 3142 4286
rect 3130 4276 3132 4284
rect 3140 4276 3142 4284
rect 2778 4124 2838 4126
rect 2778 4116 2828 4124
rect 2836 4116 2838 4124
rect 2778 4114 2838 4116
rect 2778 4104 2790 4114
rect 2778 4096 2780 4104
rect 2788 4096 2790 4104
rect 2778 4094 2790 4096
rect 2842 4084 2854 4086
rect 2842 4076 2844 4084
rect 2852 4076 2854 4084
rect 2490 4056 2492 4064
rect 2500 4056 2502 4064
rect 2490 4054 2502 4056
rect 2682 4064 2694 4066
rect 2682 4056 2684 4064
rect 2692 4056 2694 4064
rect 2458 3144 2470 3146
rect 2458 3136 2460 3144
rect 2468 3136 2470 3144
rect 2458 2924 2470 3136
rect 2458 2916 2460 2924
rect 2468 2916 2470 2924
rect 2458 2914 2470 2916
rect 2138 2676 2140 2684
rect 2148 2676 2150 2684
rect 2138 2674 2150 2676
rect 2522 2704 2534 2706
rect 2522 2696 2524 2704
rect 2532 2696 2534 2704
rect 2106 2156 2108 2164
rect 2116 2156 2118 2164
rect 2106 2154 2118 2156
rect 2426 2284 2438 2286
rect 2426 2276 2428 2284
rect 2436 2276 2438 2284
rect 1818 2116 1820 2124
rect 1828 2116 1830 2124
rect 1818 2114 1830 2116
rect 1736 2006 1740 2014
rect 1748 2006 1756 2014
rect 1764 2006 1772 2014
rect 1780 2006 1784 2014
rect 218 1964 230 1966
rect 218 1956 220 1964
rect 228 1956 230 1964
rect 218 1924 230 1956
rect 218 1916 220 1924
rect 228 1916 230 1924
rect 218 1914 230 1916
rect 1370 1924 1382 1926
rect 1370 1916 1372 1924
rect 1380 1916 1382 1924
rect 1178 1784 1190 1786
rect 1178 1776 1180 1784
rect 1188 1776 1190 1784
rect 698 1624 710 1626
rect 698 1616 700 1624
rect 708 1616 710 1624
rect 698 1484 710 1616
rect 698 1476 700 1484
rect 708 1476 710 1484
rect 698 1474 710 1476
rect 602 1184 614 1186
rect 602 1176 604 1184
rect 612 1176 614 1184
rect 410 1104 422 1106
rect 410 1096 412 1104
rect 420 1096 422 1104
rect 346 944 358 946
rect 346 936 348 944
rect 356 936 358 944
rect 186 544 198 546
rect 186 536 188 544
rect 196 536 198 544
rect 186 224 198 536
rect 346 504 358 936
rect 346 496 348 504
rect 356 496 358 504
rect 346 494 358 496
rect 410 464 422 1096
rect 602 784 614 1176
rect 602 776 604 784
rect 612 776 614 784
rect 602 774 614 776
rect 634 1084 646 1086
rect 634 1076 636 1084
rect 644 1076 646 1084
rect 634 564 646 1076
rect 1178 1084 1190 1776
rect 1178 1076 1180 1084
rect 1188 1076 1190 1084
rect 1178 1074 1190 1076
rect 1370 1104 1382 1916
rect 1370 1096 1372 1104
rect 1380 1096 1382 1104
rect 1210 924 1222 926
rect 1210 916 1212 924
rect 1220 916 1222 924
rect 1210 624 1222 916
rect 1370 864 1382 1096
rect 1736 1614 1784 2006
rect 2106 1784 2118 1786
rect 2106 1776 2108 1784
rect 2116 1776 2118 1784
rect 1736 1606 1740 1614
rect 1748 1606 1756 1614
rect 1764 1606 1772 1614
rect 1780 1606 1784 1614
rect 1736 1214 1784 1606
rect 1736 1206 1740 1214
rect 1748 1206 1756 1214
rect 1764 1206 1772 1214
rect 1780 1206 1784 1214
rect 1402 1024 1414 1026
rect 1402 1016 1404 1024
rect 1412 1016 1414 1024
rect 1402 924 1414 1016
rect 1402 916 1404 924
rect 1412 916 1414 924
rect 1402 914 1414 916
rect 1434 1004 1446 1006
rect 1434 996 1436 1004
rect 1444 996 1446 1004
rect 1434 924 1446 996
rect 1434 916 1436 924
rect 1444 916 1446 924
rect 1434 914 1446 916
rect 1530 1004 1542 1006
rect 1530 996 1532 1004
rect 1540 996 1542 1004
rect 1370 856 1372 864
rect 1380 856 1382 864
rect 1370 854 1382 856
rect 1530 704 1542 996
rect 1530 696 1532 704
rect 1540 696 1542 704
rect 1530 694 1542 696
rect 1594 904 1606 906
rect 1594 896 1596 904
rect 1604 896 1606 904
rect 1210 616 1212 624
rect 1220 616 1222 624
rect 1210 584 1222 616
rect 1594 624 1606 896
rect 1594 616 1596 624
rect 1604 616 1606 624
rect 1594 614 1606 616
rect 1736 814 1784 1206
rect 2042 1744 2054 1746
rect 2042 1736 2044 1744
rect 2052 1736 2054 1744
rect 2042 1064 2054 1736
rect 2106 1104 2118 1776
rect 2106 1096 2108 1104
rect 2116 1096 2118 1104
rect 2106 1094 2118 1096
rect 2298 1524 2310 1526
rect 2298 1516 2300 1524
rect 2308 1516 2310 1524
rect 2042 1056 2044 1064
rect 2052 1056 2054 1064
rect 2042 1054 2054 1056
rect 1736 806 1740 814
rect 1748 806 1756 814
rect 1764 806 1772 814
rect 1780 806 1784 814
rect 1210 576 1212 584
rect 1220 576 1222 584
rect 1210 574 1222 576
rect 634 556 636 564
rect 644 556 646 564
rect 634 554 646 556
rect 410 456 412 464
rect 420 456 422 464
rect 410 454 422 456
rect 186 216 188 224
rect 196 216 198 224
rect 186 214 198 216
rect 1736 414 1784 806
rect 2298 464 2310 1516
rect 2426 1364 2438 2276
rect 2522 1644 2534 2696
rect 2682 2704 2694 4056
rect 2842 4024 2854 4076
rect 2842 4016 2844 4024
rect 2852 4016 2854 4024
rect 2842 4014 2854 4016
rect 2714 4004 2726 4006
rect 2714 3996 2716 4004
rect 2724 3996 2726 4004
rect 2714 3504 2726 3996
rect 2714 3496 2716 3504
rect 2724 3496 2726 3504
rect 2714 3494 2726 3496
rect 3098 3344 3110 3346
rect 3098 3336 3100 3344
rect 3108 3336 3110 3344
rect 2810 3244 2822 3246
rect 2810 3236 2812 3244
rect 2820 3236 2822 3244
rect 2810 2844 2822 3236
rect 2810 2836 2812 2844
rect 2820 2836 2822 2844
rect 2810 2834 2822 2836
rect 3034 3064 3046 3066
rect 3034 3056 3036 3064
rect 3044 3056 3046 3064
rect 2682 2696 2684 2704
rect 2692 2696 2694 2704
rect 2682 2694 2694 2696
rect 2778 2304 2790 2306
rect 2778 2296 2780 2304
rect 2788 2296 2790 2304
rect 2746 2284 2758 2286
rect 2746 2276 2748 2284
rect 2756 2276 2758 2284
rect 2522 1636 2524 1644
rect 2532 1636 2534 1644
rect 2522 1634 2534 1636
rect 2554 2264 2566 2266
rect 2554 2256 2556 2264
rect 2564 2256 2566 2264
rect 2426 1356 2428 1364
rect 2436 1356 2438 1364
rect 2426 1354 2438 1356
rect 2554 1024 2566 2256
rect 2714 2264 2726 2266
rect 2714 2256 2716 2264
rect 2724 2256 2726 2264
rect 2714 2164 2726 2256
rect 2714 2156 2716 2164
rect 2724 2156 2726 2164
rect 2714 2154 2726 2156
rect 2746 2124 2758 2276
rect 2778 2184 2790 2296
rect 3034 2284 3046 3056
rect 3098 2684 3110 3336
rect 3130 2804 3142 4276
rect 3130 2796 3132 2804
rect 3140 2796 3142 2804
rect 3130 2794 3142 2796
rect 3162 4244 3174 4396
rect 3162 4236 3164 4244
rect 3172 4236 3174 4244
rect 3162 2864 3174 4236
rect 3272 4214 3320 4606
rect 3354 4864 3366 4866
rect 3354 4856 3356 4864
rect 3364 4856 3366 4864
rect 3354 4424 3366 4856
rect 4090 4624 4102 5236
rect 4090 4616 4092 4624
rect 4100 4616 4102 4624
rect 4090 4614 4102 4616
rect 4186 5044 4198 5046
rect 4186 5036 4188 5044
rect 4196 5036 4198 5044
rect 3354 4416 3356 4424
rect 3364 4416 3366 4424
rect 3354 4414 3366 4416
rect 3866 4584 3878 4586
rect 3866 4576 3868 4584
rect 3876 4576 3878 4584
rect 3866 4344 3878 4576
rect 3866 4336 3868 4344
rect 3876 4336 3878 4344
rect 3866 4334 3878 4336
rect 3272 4206 3276 4214
rect 3284 4206 3292 4214
rect 3300 4206 3308 4214
rect 3316 4206 3320 4214
rect 3272 3814 3320 4206
rect 3482 4304 3494 4306
rect 3482 4296 3484 4304
rect 3492 4296 3494 4304
rect 3272 3806 3276 3814
rect 3284 3806 3292 3814
rect 3300 3806 3308 3814
rect 3316 3806 3320 3814
rect 3272 3414 3320 3806
rect 3386 4184 3398 4186
rect 3386 4176 3388 4184
rect 3396 4176 3398 4184
rect 3272 3406 3276 3414
rect 3284 3406 3292 3414
rect 3300 3406 3308 3414
rect 3316 3406 3320 3414
rect 3272 3014 3320 3406
rect 3354 3484 3366 3486
rect 3354 3476 3356 3484
rect 3364 3476 3366 3484
rect 3354 3404 3366 3476
rect 3354 3396 3356 3404
rect 3364 3396 3366 3404
rect 3354 3394 3366 3396
rect 3272 3006 3276 3014
rect 3284 3006 3292 3014
rect 3300 3006 3308 3014
rect 3316 3006 3320 3014
rect 3162 2856 3164 2864
rect 3172 2856 3174 2864
rect 3098 2676 3100 2684
rect 3108 2676 3110 2684
rect 3098 2604 3110 2676
rect 3098 2596 3100 2604
rect 3108 2596 3110 2604
rect 3098 2594 3110 2596
rect 3162 2384 3174 2856
rect 3162 2376 3164 2384
rect 3172 2376 3174 2384
rect 3162 2374 3174 2376
rect 3194 2924 3206 2926
rect 3194 2916 3196 2924
rect 3204 2916 3206 2924
rect 3034 2276 3036 2284
rect 3044 2276 3046 2284
rect 3034 2274 3046 2276
rect 3066 2324 3078 2326
rect 3066 2316 3068 2324
rect 3076 2316 3078 2324
rect 2778 2176 2780 2184
rect 2788 2176 2790 2184
rect 2778 2174 2790 2176
rect 2746 2116 2748 2124
rect 2756 2116 2758 2124
rect 2746 2114 2758 2116
rect 2778 2104 2790 2106
rect 2778 2096 2780 2104
rect 2788 2096 2790 2104
rect 2778 1824 2790 2096
rect 2778 1816 2780 1824
rect 2788 1816 2790 1824
rect 2778 1814 2790 1816
rect 2842 1964 2854 1966
rect 2842 1956 2844 1964
rect 2852 1956 2854 1964
rect 2842 1744 2854 1956
rect 2874 1844 2886 1846
rect 2874 1836 2876 1844
rect 2884 1836 2886 1844
rect 2874 1764 2886 1836
rect 2874 1756 2876 1764
rect 2884 1756 2886 1764
rect 2874 1754 2886 1756
rect 2842 1736 2844 1744
rect 2852 1736 2854 1744
rect 2842 1734 2854 1736
rect 3002 1584 3014 1586
rect 3002 1576 3004 1584
rect 3012 1576 3014 1584
rect 2554 1016 2556 1024
rect 2564 1016 2566 1024
rect 2554 1014 2566 1016
rect 2650 1304 2662 1306
rect 2650 1296 2652 1304
rect 2660 1296 2662 1304
rect 2650 584 2662 1296
rect 2682 1084 2694 1086
rect 2682 1076 2684 1084
rect 2692 1076 2694 1084
rect 2682 824 2694 1076
rect 3002 1004 3014 1576
rect 3066 1504 3078 2316
rect 3066 1496 3068 1504
rect 3076 1496 3078 1504
rect 3066 1494 3078 1496
rect 3098 2004 3110 2006
rect 3098 1996 3100 2004
rect 3108 1996 3110 2004
rect 3098 1024 3110 1996
rect 3194 2004 3206 2916
rect 3194 1996 3196 2004
rect 3204 1996 3206 2004
rect 3194 1994 3206 1996
rect 3272 2614 3320 3006
rect 3386 2924 3398 4176
rect 3482 4084 3494 4296
rect 4186 4204 4198 5036
rect 4314 4524 4326 5356
rect 4730 5424 4742 5426
rect 4730 5416 4732 5424
rect 4740 5416 4742 5424
rect 4730 5324 4742 5416
rect 4730 5316 4732 5324
rect 4740 5316 4742 5324
rect 4730 5004 4742 5316
rect 4730 4996 4732 5004
rect 4740 4996 4742 5004
rect 4730 4994 4742 4996
rect 4808 5214 4856 5606
rect 5562 5564 5574 5566
rect 5562 5556 5564 5564
rect 5572 5556 5574 5564
rect 5562 5344 5574 5556
rect 5882 5504 5894 5676
rect 5882 5496 5884 5504
rect 5892 5496 5894 5504
rect 5882 5494 5894 5496
rect 5562 5336 5564 5344
rect 5572 5336 5574 5344
rect 5562 5334 5574 5336
rect 6106 5344 6118 5756
rect 6106 5336 6108 5344
rect 6116 5336 6118 5344
rect 6106 5334 6118 5336
rect 4808 5206 4812 5214
rect 4820 5206 4828 5214
rect 4836 5206 4844 5214
rect 4852 5206 4856 5214
rect 4442 4824 4454 4826
rect 4442 4816 4444 4824
rect 4452 4816 4454 4824
rect 4442 4624 4454 4816
rect 4442 4616 4444 4624
rect 4452 4616 4454 4624
rect 4442 4614 4454 4616
rect 4808 4814 4856 5206
rect 5498 5084 5510 5086
rect 5498 5076 5500 5084
rect 5508 5076 5510 5084
rect 5210 4924 5222 4926
rect 5210 4916 5212 4924
rect 5220 4916 5222 4924
rect 4808 4806 4812 4814
rect 4820 4806 4828 4814
rect 4836 4806 4844 4814
rect 4852 4806 4856 4814
rect 4314 4516 4316 4524
rect 4324 4516 4326 4524
rect 4314 4514 4326 4516
rect 4570 4604 4582 4606
rect 4570 4596 4572 4604
rect 4580 4596 4582 4604
rect 4570 4324 4582 4596
rect 4570 4316 4572 4324
rect 4580 4316 4582 4324
rect 4570 4314 4582 4316
rect 4602 4524 4614 4526
rect 4602 4516 4604 4524
rect 4612 4516 4614 4524
rect 4186 4196 4188 4204
rect 4196 4196 4198 4204
rect 4186 4194 4198 4196
rect 4506 4264 4518 4266
rect 4506 4256 4508 4264
rect 4516 4256 4518 4264
rect 4506 4204 4518 4256
rect 4506 4196 4508 4204
rect 4516 4196 4518 4204
rect 4506 4194 4518 4196
rect 3770 4184 3782 4186
rect 3770 4176 3772 4184
rect 3780 4176 3782 4184
rect 3482 4076 3484 4084
rect 3492 4076 3494 4084
rect 3482 4074 3494 4076
rect 3642 4164 3654 4166
rect 3642 4156 3644 4164
rect 3652 4156 3654 4164
rect 3482 3984 3494 3986
rect 3482 3976 3484 3984
rect 3492 3976 3494 3984
rect 3482 3884 3494 3976
rect 3610 3924 3622 3926
rect 3610 3916 3612 3924
rect 3620 3916 3622 3924
rect 3482 3876 3484 3884
rect 3492 3876 3494 3884
rect 3482 3874 3494 3876
rect 3546 3884 3558 3886
rect 3546 3876 3548 3884
rect 3556 3876 3558 3884
rect 3546 3824 3558 3876
rect 3610 3864 3622 3916
rect 3610 3856 3612 3864
rect 3620 3856 3622 3864
rect 3610 3854 3622 3856
rect 3546 3816 3548 3824
rect 3556 3816 3558 3824
rect 3546 3814 3558 3816
rect 3610 3384 3622 3386
rect 3610 3376 3612 3384
rect 3620 3376 3622 3384
rect 3610 3284 3622 3376
rect 3610 3276 3612 3284
rect 3620 3276 3622 3284
rect 3610 3274 3622 3276
rect 3642 3124 3654 4156
rect 3770 4144 3782 4176
rect 3770 4136 3772 4144
rect 3780 4136 3782 4144
rect 3770 4134 3782 4136
rect 3674 4124 3686 4126
rect 3674 4116 3676 4124
rect 3684 4116 3686 4124
rect 3674 4044 3686 4116
rect 3674 4036 3676 4044
rect 3684 4036 3686 4044
rect 3674 4034 3686 4036
rect 4538 4124 4550 4126
rect 4538 4116 4540 4124
rect 4548 4116 4550 4124
rect 3770 4004 3782 4006
rect 3770 3996 3772 4004
rect 3780 3996 3782 4004
rect 3706 3884 3718 3886
rect 3706 3876 3708 3884
rect 3716 3876 3718 3884
rect 3706 3684 3718 3876
rect 3738 3864 3750 3866
rect 3738 3856 3740 3864
rect 3748 3856 3750 3864
rect 3738 3784 3750 3856
rect 3738 3776 3740 3784
rect 3748 3776 3750 3784
rect 3738 3774 3750 3776
rect 3706 3676 3708 3684
rect 3716 3676 3718 3684
rect 3706 3674 3718 3676
rect 3642 3116 3644 3124
rect 3652 3116 3654 3124
rect 3642 2964 3654 3116
rect 3642 2956 3644 2964
rect 3652 2956 3654 2964
rect 3642 2954 3654 2956
rect 3674 3444 3686 3446
rect 3674 3436 3676 3444
rect 3684 3436 3686 3444
rect 3674 3344 3686 3436
rect 3674 3336 3676 3344
rect 3684 3336 3686 3344
rect 3386 2916 3388 2924
rect 3396 2916 3398 2924
rect 3386 2914 3398 2916
rect 3642 2924 3654 2926
rect 3642 2916 3644 2924
rect 3652 2916 3654 2924
rect 3272 2606 3276 2614
rect 3284 2606 3292 2614
rect 3300 2606 3308 2614
rect 3316 2606 3320 2614
rect 3272 2214 3320 2606
rect 3642 2504 3654 2916
rect 3674 2844 3686 3336
rect 3770 3204 3782 3996
rect 4538 3824 4550 4116
rect 4538 3816 4540 3824
rect 4548 3816 4550 3824
rect 4538 3814 4550 3816
rect 4410 3784 4422 3786
rect 4410 3776 4412 3784
rect 4420 3776 4422 3784
rect 3770 3196 3772 3204
rect 3780 3196 3782 3204
rect 3770 3194 3782 3196
rect 3930 3664 3942 3666
rect 3930 3656 3932 3664
rect 3940 3656 3942 3664
rect 3674 2836 3676 2844
rect 3684 2836 3686 2844
rect 3674 2834 3686 2836
rect 3642 2496 3644 2504
rect 3652 2496 3654 2504
rect 3642 2494 3654 2496
rect 3272 2206 3276 2214
rect 3284 2206 3292 2214
rect 3300 2206 3308 2214
rect 3316 2206 3320 2214
rect 3098 1016 3100 1024
rect 3108 1016 3110 1024
rect 3098 1014 3110 1016
rect 3272 1814 3320 2206
rect 3354 2384 3366 2386
rect 3354 2376 3356 2384
rect 3364 2376 3366 2384
rect 3354 1824 3366 2376
rect 3386 2264 3398 2266
rect 3386 2256 3388 2264
rect 3396 2256 3398 2264
rect 3386 1964 3398 2256
rect 3930 2204 3942 3656
rect 3962 3564 3974 3566
rect 3962 3556 3964 3564
rect 3972 3556 3974 3564
rect 3962 2324 3974 3556
rect 4282 3324 4294 3326
rect 4282 3316 4284 3324
rect 4292 3316 4294 3324
rect 4058 3184 4070 3186
rect 4058 3176 4060 3184
rect 4068 3176 4070 3184
rect 4058 3044 4070 3176
rect 4058 3036 4060 3044
rect 4068 3036 4070 3044
rect 4058 2384 4070 3036
rect 4218 2604 4230 2606
rect 4218 2596 4220 2604
rect 4228 2596 4230 2604
rect 4058 2376 4060 2384
rect 4068 2376 4070 2384
rect 4058 2374 4070 2376
rect 4186 2564 4198 2566
rect 4186 2556 4188 2564
rect 4196 2556 4198 2564
rect 3962 2316 3964 2324
rect 3972 2316 3974 2324
rect 3962 2314 3974 2316
rect 3994 2364 4006 2366
rect 3994 2356 3996 2364
rect 4004 2356 4006 2364
rect 3930 2196 3932 2204
rect 3940 2196 3942 2204
rect 3930 2194 3942 2196
rect 3994 2064 4006 2356
rect 4186 2284 4198 2556
rect 4218 2564 4230 2596
rect 4218 2556 4220 2564
rect 4228 2556 4230 2564
rect 4218 2554 4230 2556
rect 4250 2604 4262 2606
rect 4250 2596 4252 2604
rect 4260 2596 4262 2604
rect 4250 2304 4262 2596
rect 4282 2464 4294 3316
rect 4410 3084 4422 3776
rect 4570 3764 4582 3766
rect 4570 3756 4572 3764
rect 4580 3756 4582 3764
rect 4570 3704 4582 3756
rect 4570 3696 4572 3704
rect 4580 3696 4582 3704
rect 4570 3694 4582 3696
rect 4538 3544 4550 3546
rect 4538 3536 4540 3544
rect 4548 3536 4550 3544
rect 4538 3484 4550 3536
rect 4538 3476 4540 3484
rect 4548 3476 4550 3484
rect 4538 3474 4550 3476
rect 4410 3076 4412 3084
rect 4420 3076 4422 3084
rect 4410 3074 4422 3076
rect 4538 3044 4550 3046
rect 4538 3036 4540 3044
rect 4548 3036 4550 3044
rect 4538 2664 4550 3036
rect 4538 2656 4540 2664
rect 4548 2656 4550 2664
rect 4538 2654 4550 2656
rect 4602 2544 4614 4516
rect 4808 4414 4856 4806
rect 5050 4844 5062 4846
rect 5050 4836 5052 4844
rect 5060 4836 5062 4844
rect 5050 4624 5062 4836
rect 5050 4616 5052 4624
rect 5060 4616 5062 4624
rect 5050 4424 5062 4616
rect 5050 4416 5052 4424
rect 5060 4416 5062 4424
rect 5050 4414 5062 4416
rect 5178 4464 5190 4466
rect 5178 4456 5180 4464
rect 5188 4456 5190 4464
rect 4808 4406 4812 4414
rect 4820 4406 4828 4414
rect 4836 4406 4844 4414
rect 4852 4406 4856 4414
rect 4730 4244 4742 4246
rect 4730 4236 4732 4244
rect 4740 4236 4742 4244
rect 4698 3644 4710 3646
rect 4698 3636 4700 3644
rect 4708 3636 4710 3644
rect 4634 3604 4646 3606
rect 4634 3596 4636 3604
rect 4644 3596 4646 3604
rect 4634 3344 4646 3596
rect 4634 3336 4636 3344
rect 4644 3336 4646 3344
rect 4634 3334 4646 3336
rect 4666 3064 4678 3066
rect 4666 3056 4668 3064
rect 4676 3056 4678 3064
rect 4602 2536 4604 2544
rect 4612 2536 4614 2544
rect 4602 2534 4614 2536
rect 4634 2804 4646 2806
rect 4634 2796 4636 2804
rect 4644 2796 4646 2804
rect 4282 2456 4284 2464
rect 4292 2456 4294 2464
rect 4282 2454 4294 2456
rect 4250 2296 4252 2304
rect 4260 2296 4262 2304
rect 4250 2294 4262 2296
rect 4314 2424 4326 2426
rect 4314 2416 4316 2424
rect 4324 2416 4326 2424
rect 4186 2276 4188 2284
rect 4196 2276 4198 2284
rect 4186 2144 4198 2276
rect 4186 2136 4188 2144
rect 4196 2136 4198 2144
rect 4186 2134 4198 2136
rect 4314 2144 4326 2416
rect 4314 2136 4316 2144
rect 4324 2136 4326 2144
rect 4314 2134 4326 2136
rect 4410 2424 4422 2426
rect 4410 2416 4412 2424
rect 4420 2416 4422 2424
rect 3994 2056 3996 2064
rect 4004 2056 4006 2064
rect 3994 2054 4006 2056
rect 3386 1956 3388 1964
rect 3396 1956 3398 1964
rect 3386 1954 3398 1956
rect 4410 1904 4422 2416
rect 4410 1896 4412 1904
rect 4420 1896 4422 1904
rect 4410 1894 4422 1896
rect 4538 2024 4550 2026
rect 4538 2016 4540 2024
rect 4548 2016 4550 2024
rect 3354 1816 3356 1824
rect 3364 1816 3366 1824
rect 3354 1814 3366 1816
rect 3962 1884 3974 1886
rect 3962 1876 3964 1884
rect 3972 1876 3974 1884
rect 3272 1806 3276 1814
rect 3284 1806 3292 1814
rect 3300 1806 3308 1814
rect 3316 1806 3320 1814
rect 3272 1414 3320 1806
rect 3770 1784 3782 1786
rect 3770 1776 3772 1784
rect 3780 1776 3782 1784
rect 3418 1744 3430 1746
rect 3418 1736 3420 1744
rect 3428 1736 3430 1744
rect 3418 1684 3430 1736
rect 3770 1704 3782 1776
rect 3770 1696 3772 1704
rect 3780 1696 3782 1704
rect 3770 1694 3782 1696
rect 3418 1676 3420 1684
rect 3428 1676 3430 1684
rect 3418 1674 3430 1676
rect 3272 1406 3276 1414
rect 3284 1406 3292 1414
rect 3300 1406 3308 1414
rect 3316 1406 3320 1414
rect 3272 1014 3320 1406
rect 3450 1504 3462 1506
rect 3450 1496 3452 1504
rect 3460 1496 3462 1504
rect 3002 996 3004 1004
rect 3012 996 3014 1004
rect 3002 994 3014 996
rect 3272 1006 3276 1014
rect 3284 1006 3292 1014
rect 3300 1006 3308 1014
rect 3316 1006 3320 1014
rect 2682 816 2684 824
rect 2692 816 2694 824
rect 2682 814 2694 816
rect 2650 576 2652 584
rect 2660 576 2662 584
rect 2650 574 2662 576
rect 3272 614 3320 1006
rect 3272 606 3276 614
rect 3284 606 3292 614
rect 3300 606 3308 614
rect 3316 606 3320 614
rect 2298 456 2300 464
rect 2308 456 2310 464
rect 2298 454 2310 456
rect 1736 406 1740 414
rect 1748 406 1756 414
rect 1764 406 1772 414
rect 1780 406 1784 414
rect 1736 14 1784 406
rect 3226 384 3238 386
rect 3226 376 3228 384
rect 3236 376 3238 384
rect 2714 324 2726 326
rect 2714 316 2716 324
rect 2724 316 2726 324
rect 2714 284 2726 316
rect 2714 276 2716 284
rect 2724 276 2726 284
rect 2714 274 2726 276
rect 2074 184 2086 186
rect 2074 176 2076 184
rect 2084 176 2086 184
rect 2074 166 2086 176
rect 2074 164 2150 166
rect 2074 156 2140 164
rect 2148 156 2150 164
rect 2074 154 2150 156
rect 3226 144 3238 376
rect 3226 136 3228 144
rect 3236 136 3238 144
rect 3226 134 3238 136
rect 3272 214 3320 606
rect 3354 1204 3366 1206
rect 3354 1196 3356 1204
rect 3364 1196 3366 1204
rect 3354 444 3366 1196
rect 3450 664 3462 1496
rect 3706 1104 3718 1106
rect 3706 1096 3708 1104
rect 3716 1096 3718 1104
rect 3674 1064 3686 1066
rect 3674 1056 3676 1064
rect 3684 1056 3686 1064
rect 3674 944 3686 1056
rect 3674 936 3676 944
rect 3684 936 3686 944
rect 3674 934 3686 936
rect 3706 744 3718 1096
rect 3706 736 3708 744
rect 3716 736 3718 744
rect 3706 704 3718 736
rect 3866 1104 3878 1106
rect 3866 1096 3868 1104
rect 3876 1096 3878 1104
rect 3866 724 3878 1096
rect 3930 1064 3942 1066
rect 3930 1056 3932 1064
rect 3940 1056 3942 1064
rect 3930 1024 3942 1056
rect 3930 1016 3932 1024
rect 3940 1016 3942 1024
rect 3930 1014 3942 1016
rect 3866 716 3868 724
rect 3876 716 3878 724
rect 3866 714 3878 716
rect 3706 696 3708 704
rect 3716 696 3718 704
rect 3706 694 3718 696
rect 3450 656 3452 664
rect 3460 656 3462 664
rect 3450 654 3462 656
rect 3962 664 3974 1876
rect 4474 1764 4486 1766
rect 4474 1756 4476 1764
rect 4484 1756 4486 1764
rect 4410 1744 4422 1746
rect 4410 1736 4412 1744
rect 4420 1736 4422 1744
rect 4090 1724 4102 1726
rect 4090 1716 4092 1724
rect 4100 1716 4102 1724
rect 4090 1424 4102 1716
rect 4090 1416 4092 1424
rect 4100 1416 4102 1424
rect 4090 1414 4102 1416
rect 4378 1664 4390 1666
rect 4378 1656 4380 1664
rect 4388 1656 4390 1664
rect 4250 1184 4262 1186
rect 4250 1176 4252 1184
rect 4260 1176 4262 1184
rect 4250 764 4262 1176
rect 4346 1064 4358 1066
rect 4346 1056 4348 1064
rect 4356 1056 4358 1064
rect 4346 1004 4358 1056
rect 4346 996 4348 1004
rect 4356 996 4358 1004
rect 4346 924 4358 996
rect 4346 916 4348 924
rect 4356 916 4358 924
rect 4346 914 4358 916
rect 4250 756 4252 764
rect 4260 756 4262 764
rect 4250 754 4262 756
rect 4378 684 4390 1656
rect 4410 1664 4422 1736
rect 4410 1656 4412 1664
rect 4420 1656 4422 1664
rect 4410 1654 4422 1656
rect 4378 676 4380 684
rect 4388 676 4390 684
rect 4378 674 4390 676
rect 4474 784 4486 1756
rect 4506 1704 4518 1706
rect 4506 1696 4508 1704
rect 4516 1696 4518 1704
rect 4506 1624 4518 1696
rect 4506 1616 4508 1624
rect 4516 1616 4518 1624
rect 4506 1614 4518 1616
rect 4538 1424 4550 2016
rect 4634 2024 4646 2796
rect 4666 2684 4678 3056
rect 4698 2804 4710 3636
rect 4730 3644 4742 4236
rect 4730 3636 4732 3644
rect 4740 3636 4742 3644
rect 4730 3634 4742 3636
rect 4808 4014 4856 4406
rect 4986 4304 4998 4306
rect 4986 4296 4988 4304
rect 4996 4296 4998 4304
rect 4808 4006 4812 4014
rect 4820 4006 4828 4014
rect 4836 4006 4844 4014
rect 4852 4006 4856 4014
rect 4698 2796 4700 2804
rect 4708 2796 4710 2804
rect 4698 2794 4710 2796
rect 4808 3614 4856 4006
rect 4890 4144 4902 4146
rect 4890 4136 4892 4144
rect 4900 4136 4902 4144
rect 4890 3824 4902 4136
rect 4986 4124 4998 4296
rect 4986 4116 4988 4124
rect 4996 4116 4998 4124
rect 4986 4114 4998 4116
rect 5050 4284 5062 4286
rect 5050 4276 5052 4284
rect 5060 4276 5062 4284
rect 4890 3816 4892 3824
rect 4900 3816 4902 3824
rect 4890 3814 4902 3816
rect 5050 4024 5062 4276
rect 5178 4064 5190 4456
rect 5178 4056 5180 4064
rect 5188 4056 5190 4064
rect 5178 4054 5190 4056
rect 5050 4016 5052 4024
rect 5060 4016 5062 4024
rect 4808 3606 4812 3614
rect 4820 3606 4828 3614
rect 4836 3606 4844 3614
rect 4852 3606 4856 3614
rect 4808 3214 4856 3606
rect 4808 3206 4812 3214
rect 4820 3206 4828 3214
rect 4836 3206 4844 3214
rect 4852 3206 4856 3214
rect 4808 2814 4856 3206
rect 4922 3664 4934 3666
rect 4922 3656 4924 3664
rect 4932 3656 4934 3664
rect 4890 3184 4902 3186
rect 4890 3176 4892 3184
rect 4900 3176 4902 3184
rect 4890 2904 4902 3176
rect 4890 2896 4892 2904
rect 4900 2896 4902 2904
rect 4890 2894 4902 2896
rect 4808 2806 4812 2814
rect 4820 2806 4828 2814
rect 4836 2806 4844 2814
rect 4852 2806 4856 2814
rect 4666 2676 4668 2684
rect 4676 2676 4678 2684
rect 4666 2164 4678 2676
rect 4698 2484 4710 2486
rect 4698 2476 4700 2484
rect 4708 2476 4710 2484
rect 4698 2184 4710 2476
rect 4808 2414 4856 2806
rect 4808 2406 4812 2414
rect 4820 2406 4828 2414
rect 4836 2406 4844 2414
rect 4852 2406 4856 2414
rect 4762 2364 4774 2366
rect 4762 2356 4764 2364
rect 4772 2356 4774 2364
rect 4762 2324 4774 2356
rect 4762 2316 4764 2324
rect 4772 2316 4774 2324
rect 4762 2314 4774 2316
rect 4698 2176 4700 2184
rect 4708 2176 4710 2184
rect 4698 2174 4710 2176
rect 4666 2156 4668 2164
rect 4676 2156 4678 2164
rect 4666 2154 4678 2156
rect 4634 2016 4636 2024
rect 4644 2016 4646 2024
rect 4634 2014 4646 2016
rect 4808 2014 4856 2406
rect 4808 2006 4812 2014
rect 4820 2006 4828 2014
rect 4836 2006 4844 2014
rect 4852 2006 4856 2014
rect 4602 1904 4614 1906
rect 4602 1896 4604 1904
rect 4612 1896 4614 1904
rect 4602 1804 4614 1896
rect 4602 1796 4604 1804
rect 4612 1796 4614 1804
rect 4602 1794 4614 1796
rect 4538 1416 4540 1424
rect 4548 1416 4550 1424
rect 4538 1414 4550 1416
rect 4808 1614 4856 2006
rect 4808 1606 4812 1614
rect 4820 1606 4828 1614
rect 4836 1606 4844 1614
rect 4852 1606 4856 1614
rect 4474 776 4476 784
rect 4484 776 4486 784
rect 3962 656 3964 664
rect 3972 656 3974 664
rect 3962 654 3974 656
rect 3354 436 3356 444
rect 3364 436 3366 444
rect 3354 434 3366 436
rect 3578 484 3590 486
rect 3578 476 3580 484
rect 3588 476 3590 484
rect 3578 244 3590 476
rect 4474 444 4486 776
rect 4808 1214 4856 1606
rect 4922 1284 4934 3656
rect 4986 3644 4998 3646
rect 4986 3636 4988 3644
rect 4996 3636 4998 3644
rect 4986 2444 4998 3636
rect 5050 2844 5062 4016
rect 5146 3504 5158 3506
rect 5146 3496 5148 3504
rect 5156 3496 5158 3504
rect 5146 3404 5158 3496
rect 5146 3396 5148 3404
rect 5156 3396 5158 3404
rect 5146 3394 5158 3396
rect 5082 3324 5094 3326
rect 5082 3316 5084 3324
rect 5092 3316 5094 3324
rect 5082 3284 5094 3316
rect 5210 3304 5222 4916
rect 5338 4704 5350 4706
rect 5338 4696 5340 4704
rect 5348 4696 5350 4704
rect 5338 4644 5350 4696
rect 5338 4636 5340 4644
rect 5348 4636 5350 4644
rect 5338 4634 5350 4636
rect 5466 4704 5478 4706
rect 5466 4696 5468 4704
rect 5476 4696 5478 4704
rect 5402 4244 5414 4246
rect 5402 4236 5404 4244
rect 5412 4236 5414 4244
rect 5274 4184 5286 4186
rect 5274 4176 5276 4184
rect 5284 4176 5286 4184
rect 5274 4124 5286 4176
rect 5274 4116 5276 4124
rect 5284 4116 5286 4124
rect 5274 4114 5286 4116
rect 5338 4164 5350 4166
rect 5338 4156 5340 4164
rect 5348 4156 5350 4164
rect 5338 3604 5350 4156
rect 5338 3596 5340 3604
rect 5348 3596 5350 3604
rect 5338 3594 5350 3596
rect 5370 3604 5382 3606
rect 5370 3596 5372 3604
rect 5380 3596 5382 3604
rect 5210 3296 5212 3304
rect 5220 3296 5222 3304
rect 5210 3294 5222 3296
rect 5082 3276 5084 3284
rect 5092 3276 5094 3284
rect 5082 3274 5094 3276
rect 5050 2836 5052 2844
rect 5060 2836 5062 2844
rect 5050 2834 5062 2836
rect 5146 2924 5158 2926
rect 5146 2916 5148 2924
rect 5156 2916 5158 2924
rect 5146 2644 5158 2916
rect 5146 2636 5148 2644
rect 5156 2636 5158 2644
rect 5146 2634 5158 2636
rect 5370 2484 5382 3596
rect 5402 3544 5414 4236
rect 5402 3536 5404 3544
rect 5412 3536 5414 3544
rect 5402 3534 5414 3536
rect 5466 3784 5478 4696
rect 5466 3776 5468 3784
rect 5476 3776 5478 3784
rect 5466 3384 5478 3776
rect 5498 4004 5510 5076
rect 5562 5044 5574 5046
rect 5562 5036 5564 5044
rect 5572 5036 5574 5044
rect 5498 3996 5500 4004
rect 5508 3996 5510 4004
rect 5498 3764 5510 3996
rect 5498 3756 5500 3764
rect 5508 3756 5510 3764
rect 5498 3754 5510 3756
rect 5530 4324 5542 4326
rect 5530 4316 5532 4324
rect 5540 4316 5542 4324
rect 5530 3764 5542 4316
rect 5562 4304 5574 5036
rect 5786 4884 5798 4886
rect 5786 4876 5788 4884
rect 5796 4876 5798 4884
rect 5786 4644 5798 4876
rect 5786 4636 5788 4644
rect 5796 4636 5798 4644
rect 5786 4634 5798 4636
rect 6138 4464 6150 4466
rect 6138 4456 6140 4464
rect 6148 4456 6150 4464
rect 5562 4296 5564 4304
rect 5572 4296 5574 4304
rect 5562 4294 5574 4296
rect 5946 4444 5958 4446
rect 5946 4436 5948 4444
rect 5956 4436 5958 4444
rect 5530 3756 5532 3764
rect 5540 3756 5542 3764
rect 5530 3754 5542 3756
rect 5914 4044 5926 4046
rect 5914 4036 5916 4044
rect 5924 4036 5926 4044
rect 5466 3376 5468 3384
rect 5476 3376 5478 3384
rect 5466 3374 5478 3376
rect 5882 3624 5894 3626
rect 5882 3616 5884 3624
rect 5892 3616 5894 3624
rect 5562 2984 5574 2986
rect 5562 2976 5564 2984
rect 5572 2976 5574 2984
rect 5370 2476 5372 2484
rect 5380 2476 5382 2484
rect 5370 2474 5382 2476
rect 5434 2844 5446 2846
rect 5434 2836 5436 2844
rect 5444 2836 5446 2844
rect 4986 2436 4988 2444
rect 4996 2436 4998 2444
rect 4986 2434 4998 2436
rect 5434 1984 5446 2836
rect 5434 1976 5436 1984
rect 5444 1976 5446 1984
rect 5434 1974 5446 1976
rect 5562 2504 5574 2976
rect 5882 2804 5894 3616
rect 5882 2796 5884 2804
rect 5892 2796 5894 2804
rect 5882 2794 5894 2796
rect 5562 2496 5564 2504
rect 5572 2496 5574 2504
rect 5562 1904 5574 2496
rect 5914 2364 5926 4036
rect 5946 3904 5958 4436
rect 6138 4184 6150 4456
rect 6138 4176 6140 4184
rect 6148 4176 6150 4184
rect 6138 4174 6150 4176
rect 6202 4044 6214 5796
rect 6344 5414 6392 5806
rect 6344 5406 6348 5414
rect 6356 5406 6364 5414
rect 6372 5406 6380 5414
rect 6388 5406 6392 5414
rect 6344 5014 6392 5406
rect 7354 5744 7366 5746
rect 7354 5736 7356 5744
rect 7364 5736 7366 5744
rect 7066 5364 7078 5366
rect 7066 5356 7068 5364
rect 7076 5356 7078 5364
rect 7066 5304 7078 5356
rect 7066 5296 7068 5304
rect 7076 5296 7078 5304
rect 7066 5294 7078 5296
rect 6906 5104 6918 5106
rect 6906 5096 6908 5104
rect 6916 5096 6918 5104
rect 6906 5044 6918 5096
rect 6906 5036 6908 5044
rect 6916 5036 6918 5044
rect 6906 5034 6918 5036
rect 7162 5064 7174 5066
rect 7162 5056 7164 5064
rect 7172 5056 7174 5064
rect 6344 5006 6348 5014
rect 6356 5006 6364 5014
rect 6372 5006 6380 5014
rect 6388 5006 6392 5014
rect 6344 4614 6392 5006
rect 7162 4664 7174 5056
rect 7226 4984 7238 4986
rect 7226 4976 7228 4984
rect 7236 4976 7238 4984
rect 7226 4924 7238 4976
rect 7354 4984 7366 5736
rect 7642 5744 7654 5746
rect 7642 5736 7644 5744
rect 7652 5736 7654 5744
rect 7450 5624 7462 5626
rect 7450 5616 7452 5624
rect 7460 5616 7462 5624
rect 7354 4976 7356 4984
rect 7364 4976 7366 4984
rect 7354 4974 7366 4976
rect 7418 5584 7430 5586
rect 7418 5576 7420 5584
rect 7428 5576 7430 5584
rect 7226 4916 7228 4924
rect 7236 4916 7238 4924
rect 7226 4914 7238 4916
rect 7162 4656 7164 4664
rect 7172 4656 7174 4664
rect 7162 4654 7174 4656
rect 6344 4606 6348 4614
rect 6356 4606 6364 4614
rect 6372 4606 6380 4614
rect 6388 4606 6392 4614
rect 6298 4284 6310 4286
rect 6298 4276 6300 4284
rect 6308 4276 6310 4284
rect 6298 4124 6310 4276
rect 6298 4116 6300 4124
rect 6308 4116 6310 4124
rect 6298 4114 6310 4116
rect 6344 4214 6392 4606
rect 6344 4206 6348 4214
rect 6356 4206 6364 4214
rect 6372 4206 6380 4214
rect 6388 4206 6392 4214
rect 6202 4036 6204 4044
rect 6212 4036 6214 4044
rect 6202 4034 6214 4036
rect 5946 3896 5948 3904
rect 5956 3896 5958 3904
rect 5946 3894 5958 3896
rect 6106 4004 6118 4006
rect 6106 3996 6108 4004
rect 6116 3996 6118 4004
rect 6074 3464 6086 3466
rect 6074 3456 6076 3464
rect 6084 3456 6086 3464
rect 6074 3344 6086 3456
rect 6106 3424 6118 3996
rect 6234 3884 6246 3886
rect 6234 3876 6236 3884
rect 6244 3876 6246 3884
rect 6106 3416 6108 3424
rect 6116 3416 6118 3424
rect 6106 3414 6118 3416
rect 6138 3584 6150 3586
rect 6138 3576 6140 3584
rect 6148 3576 6150 3584
rect 6074 3336 6076 3344
rect 6084 3336 6086 3344
rect 6074 3334 6086 3336
rect 6138 2824 6150 3576
rect 6234 3184 6246 3876
rect 6344 3814 6392 4206
rect 6490 4584 6502 4586
rect 6490 4576 6492 4584
rect 6500 4576 6502 4584
rect 6490 4204 6502 4576
rect 7290 4484 7302 4486
rect 7290 4476 7292 4484
rect 7300 4476 7302 4484
rect 6490 4196 6492 4204
rect 6500 4196 6502 4204
rect 6490 4194 6502 4196
rect 6682 4284 6694 4286
rect 6682 4276 6684 4284
rect 6692 4276 6694 4284
rect 6682 4144 6694 4276
rect 6682 4136 6684 4144
rect 6692 4136 6694 4144
rect 6344 3806 6348 3814
rect 6356 3806 6364 3814
rect 6372 3806 6380 3814
rect 6388 3806 6392 3814
rect 6234 3176 6236 3184
rect 6244 3176 6246 3184
rect 6234 3174 6246 3176
rect 6266 3684 6278 3686
rect 6266 3676 6268 3684
rect 6276 3676 6278 3684
rect 6266 3084 6278 3676
rect 6266 3076 6268 3084
rect 6276 3076 6278 3084
rect 6266 3074 6278 3076
rect 6344 3414 6392 3806
rect 6618 3904 6630 3906
rect 6618 3896 6620 3904
rect 6628 3896 6630 3904
rect 6618 3804 6630 3896
rect 6618 3796 6620 3804
rect 6628 3796 6630 3804
rect 6618 3794 6630 3796
rect 6344 3406 6348 3414
rect 6356 3406 6364 3414
rect 6372 3406 6380 3414
rect 6388 3406 6392 3414
rect 6138 2816 6140 2824
rect 6148 2816 6150 2824
rect 6138 2814 6150 2816
rect 6344 3014 6392 3406
rect 6344 3006 6348 3014
rect 6356 3006 6364 3014
rect 6372 3006 6380 3014
rect 6388 3006 6392 3014
rect 6298 2744 6310 2746
rect 6298 2736 6300 2744
rect 6308 2736 6310 2744
rect 5946 2724 5958 2726
rect 5946 2716 5948 2724
rect 5956 2716 5958 2724
rect 5946 2404 5958 2716
rect 6266 2664 6278 2666
rect 6266 2656 6268 2664
rect 6276 2656 6278 2664
rect 5946 2396 5948 2404
rect 5956 2396 5958 2404
rect 5946 2394 5958 2396
rect 6202 2624 6214 2626
rect 6202 2616 6204 2624
rect 6212 2616 6214 2624
rect 5914 2356 5916 2364
rect 5924 2356 5926 2364
rect 5914 2354 5926 2356
rect 6138 2344 6150 2346
rect 6138 2336 6140 2344
rect 6148 2336 6150 2344
rect 5562 1896 5564 1904
rect 5572 1896 5574 1904
rect 5562 1894 5574 1896
rect 5690 2244 5702 2246
rect 5690 2236 5692 2244
rect 5700 2236 5702 2244
rect 5690 1904 5702 2236
rect 5690 1896 5692 1904
rect 5700 1896 5702 1904
rect 5690 1894 5702 1896
rect 5690 1824 5702 1826
rect 5690 1816 5692 1824
rect 5700 1816 5702 1824
rect 5690 1724 5702 1816
rect 6138 1784 6150 2336
rect 6202 2144 6214 2616
rect 6202 2136 6204 2144
rect 6212 2136 6214 2144
rect 6202 2134 6214 2136
rect 6234 2624 6246 2626
rect 6234 2616 6236 2624
rect 6244 2616 6246 2624
rect 6234 2144 6246 2616
rect 6266 2524 6278 2656
rect 6266 2516 6268 2524
rect 6276 2516 6278 2524
rect 6266 2514 6278 2516
rect 6298 2164 6310 2736
rect 6298 2156 6300 2164
rect 6308 2156 6310 2164
rect 6298 2154 6310 2156
rect 6344 2614 6392 3006
rect 6426 3784 6438 3786
rect 6426 3776 6428 3784
rect 6436 3776 6438 3784
rect 6426 3004 6438 3776
rect 6490 3764 6502 3766
rect 6490 3756 6492 3764
rect 6500 3756 6502 3764
rect 6490 3504 6502 3756
rect 6490 3496 6492 3504
rect 6500 3496 6502 3504
rect 6490 3494 6502 3496
rect 6618 3724 6630 3726
rect 6618 3716 6620 3724
rect 6628 3716 6630 3724
rect 6618 3644 6630 3716
rect 6618 3636 6620 3644
rect 6628 3636 6630 3644
rect 6426 2996 6428 3004
rect 6436 2996 6438 3004
rect 6426 2994 6438 2996
rect 6458 3184 6470 3186
rect 6458 3176 6460 3184
rect 6468 3176 6470 3184
rect 6344 2606 6348 2614
rect 6356 2606 6364 2614
rect 6372 2606 6380 2614
rect 6388 2606 6392 2614
rect 6344 2214 6392 2606
rect 6344 2206 6348 2214
rect 6356 2206 6364 2214
rect 6372 2206 6380 2214
rect 6388 2206 6392 2214
rect 6234 2136 6236 2144
rect 6244 2136 6246 2144
rect 6138 1776 6140 1784
rect 6148 1776 6150 1784
rect 6138 1774 6150 1776
rect 5690 1716 5692 1724
rect 5700 1716 5702 1724
rect 5690 1714 5702 1716
rect 6234 1744 6246 2136
rect 6234 1736 6236 1744
rect 6244 1736 6246 1744
rect 4922 1276 4924 1284
rect 4932 1276 4934 1284
rect 4922 1274 4934 1276
rect 5082 1584 5094 1586
rect 5082 1576 5084 1584
rect 5092 1576 5094 1584
rect 4808 1206 4812 1214
rect 4820 1206 4828 1214
rect 4836 1206 4844 1214
rect 4852 1206 4856 1214
rect 4808 814 4856 1206
rect 5082 1104 5094 1576
rect 5818 1504 5830 1506
rect 5818 1496 5820 1504
rect 5828 1496 5830 1504
rect 5818 1304 5830 1496
rect 5946 1424 5958 1426
rect 5946 1416 5948 1424
rect 5956 1416 5958 1424
rect 5818 1296 5820 1304
rect 5828 1296 5830 1304
rect 5818 1294 5830 1296
rect 5914 1364 5926 1366
rect 5914 1356 5916 1364
rect 5924 1356 5926 1364
rect 5082 1096 5084 1104
rect 5092 1096 5094 1104
rect 5082 944 5094 1096
rect 5082 936 5084 944
rect 5092 936 5094 944
rect 5082 934 5094 936
rect 5466 984 5478 986
rect 5466 976 5468 984
rect 5476 976 5478 984
rect 4808 806 4812 814
rect 4820 806 4828 814
rect 4836 806 4844 814
rect 4852 806 4856 814
rect 4698 684 4710 686
rect 4698 676 4700 684
rect 4708 676 4710 684
rect 4698 624 4710 676
rect 4698 616 4700 624
rect 4708 616 4710 624
rect 4698 614 4710 616
rect 4474 436 4476 444
rect 4484 436 4486 444
rect 4474 434 4486 436
rect 4808 414 4856 806
rect 4808 406 4812 414
rect 4820 406 4828 414
rect 4836 406 4844 414
rect 4852 406 4856 414
rect 3578 236 3580 244
rect 3588 236 3590 244
rect 3578 234 3590 236
rect 3738 284 3750 286
rect 3738 276 3740 284
rect 3748 276 3750 284
rect 3272 206 3276 214
rect 3284 206 3292 214
rect 3300 206 3308 214
rect 3316 206 3320 214
rect 1736 6 1740 14
rect 1748 6 1756 14
rect 1764 6 1772 14
rect 1780 6 1784 14
rect 1736 0 1784 6
rect 3272 0 3320 206
rect 3738 184 3750 276
rect 3738 176 3740 184
rect 3748 176 3750 184
rect 3738 174 3750 176
rect 4808 14 4856 406
rect 5466 304 5478 976
rect 5914 984 5926 1356
rect 5946 1184 5958 1416
rect 6234 1344 6246 1736
rect 6234 1336 6236 1344
rect 6244 1336 6246 1344
rect 6234 1334 6246 1336
rect 6344 1814 6392 2206
rect 6344 1806 6348 1814
rect 6356 1806 6364 1814
rect 6372 1806 6380 1814
rect 6388 1806 6392 1814
rect 6344 1414 6392 1806
rect 6426 2524 6438 2526
rect 6426 2516 6428 2524
rect 6436 2516 6438 2524
rect 6426 1504 6438 2516
rect 6458 2344 6470 3176
rect 6618 2524 6630 3636
rect 6650 3124 6662 3126
rect 6650 3116 6652 3124
rect 6660 3116 6662 3124
rect 6650 3064 6662 3116
rect 6650 3056 6652 3064
rect 6660 3056 6662 3064
rect 6650 3054 6662 3056
rect 6682 2684 6694 4136
rect 7130 4244 7142 4246
rect 7130 4236 7132 4244
rect 7140 4236 7142 4244
rect 6906 3944 6918 3946
rect 6906 3936 6908 3944
rect 6916 3936 6918 3944
rect 6906 3344 6918 3936
rect 7034 3764 7046 3766
rect 7034 3756 7036 3764
rect 7044 3756 7046 3764
rect 6906 3336 6908 3344
rect 6916 3336 6918 3344
rect 6906 3334 6918 3336
rect 6970 3564 6982 3566
rect 6970 3556 6972 3564
rect 6980 3556 6982 3564
rect 6682 2676 6684 2684
rect 6692 2676 6694 2684
rect 6682 2674 6694 2676
rect 6618 2516 6620 2524
rect 6628 2516 6630 2524
rect 6618 2514 6630 2516
rect 6458 2336 6460 2344
rect 6468 2336 6470 2344
rect 6458 2334 6470 2336
rect 6842 2364 6854 2366
rect 6842 2356 6844 2364
rect 6852 2356 6854 2364
rect 6714 2244 6726 2246
rect 6714 2236 6716 2244
rect 6724 2236 6726 2244
rect 6522 1784 6534 1786
rect 6522 1776 6524 1784
rect 6532 1776 6534 1784
rect 6522 1544 6534 1776
rect 6522 1536 6524 1544
rect 6532 1536 6534 1544
rect 6522 1534 6534 1536
rect 6714 1524 6726 2236
rect 6842 1924 6854 2356
rect 6842 1916 6844 1924
rect 6852 1916 6854 1924
rect 6842 1914 6854 1916
rect 6714 1516 6716 1524
rect 6724 1516 6726 1524
rect 6714 1514 6726 1516
rect 6426 1496 6428 1504
rect 6436 1496 6438 1504
rect 6426 1494 6438 1496
rect 6970 1504 6982 3556
rect 7034 2364 7046 3756
rect 7130 3704 7142 4236
rect 7290 3884 7302 4476
rect 7418 4424 7430 5576
rect 7418 4416 7420 4424
rect 7428 4416 7430 4424
rect 7418 4414 7430 4416
rect 7450 3944 7462 5616
rect 7610 4964 7622 4966
rect 7610 4956 7612 4964
rect 7620 4956 7622 4964
rect 7578 4724 7590 4726
rect 7578 4716 7580 4724
rect 7588 4716 7590 4724
rect 7546 4604 7558 4606
rect 7546 4596 7548 4604
rect 7556 4596 7558 4604
rect 7514 4404 7526 4406
rect 7514 4396 7516 4404
rect 7524 4396 7526 4404
rect 7514 4144 7526 4396
rect 7514 4136 7516 4144
rect 7524 4136 7526 4144
rect 7514 4134 7526 4136
rect 7450 3936 7452 3944
rect 7460 3936 7462 3944
rect 7450 3934 7462 3936
rect 7290 3876 7292 3884
rect 7300 3876 7302 3884
rect 7290 3874 7302 3876
rect 7130 3696 7132 3704
rect 7140 3696 7142 3704
rect 7130 3694 7142 3696
rect 7386 3484 7398 3486
rect 7386 3476 7388 3484
rect 7396 3476 7398 3484
rect 7290 3244 7302 3246
rect 7290 3236 7292 3244
rect 7300 3236 7302 3244
rect 7290 3084 7302 3236
rect 7290 3076 7292 3084
rect 7300 3076 7302 3084
rect 7290 2904 7302 3076
rect 7386 2964 7398 3476
rect 7546 3444 7558 4596
rect 7578 4564 7590 4716
rect 7578 4556 7580 4564
rect 7588 4556 7590 4564
rect 7578 4554 7590 4556
rect 7610 4544 7622 4956
rect 7642 4864 7654 5736
rect 7866 5744 7878 5746
rect 7866 5736 7868 5744
rect 7876 5736 7878 5744
rect 7770 5384 7782 5386
rect 7770 5376 7772 5384
rect 7780 5376 7782 5384
rect 7642 4856 7644 4864
rect 7652 4856 7654 4864
rect 7642 4854 7654 4856
rect 7674 5024 7686 5026
rect 7674 5016 7676 5024
rect 7684 5016 7686 5024
rect 7610 4536 7612 4544
rect 7620 4536 7622 4544
rect 7610 4534 7622 4536
rect 7674 4324 7686 5016
rect 7738 4944 7750 4946
rect 7738 4936 7740 4944
rect 7748 4936 7750 4944
rect 7674 4316 7676 4324
rect 7684 4316 7686 4324
rect 7674 4314 7686 4316
rect 7706 4624 7718 4626
rect 7706 4616 7708 4624
rect 7716 4616 7718 4624
rect 7706 4224 7718 4616
rect 7738 4524 7750 4936
rect 7738 4516 7740 4524
rect 7748 4516 7750 4524
rect 7738 4514 7750 4516
rect 7770 4284 7782 5376
rect 7770 4276 7772 4284
rect 7780 4276 7782 4284
rect 7770 4274 7782 4276
rect 7834 5104 7846 5106
rect 7834 5096 7836 5104
rect 7844 5096 7846 5104
rect 7706 4216 7708 4224
rect 7716 4216 7718 4224
rect 7706 4214 7718 4216
rect 7802 4084 7814 4086
rect 7802 4076 7804 4084
rect 7812 4076 7814 4084
rect 7738 4064 7750 4066
rect 7738 4056 7740 4064
rect 7748 4056 7750 4064
rect 7546 3436 7548 3444
rect 7556 3436 7558 3444
rect 7546 3434 7558 3436
rect 7674 3944 7686 3946
rect 7674 3936 7676 3944
rect 7684 3936 7686 3944
rect 7386 2956 7388 2964
rect 7396 2956 7398 2964
rect 7386 2954 7398 2956
rect 7450 3344 7462 3346
rect 7450 3336 7452 3344
rect 7460 3336 7462 3344
rect 7290 2896 7292 2904
rect 7300 2896 7302 2904
rect 7290 2894 7302 2896
rect 7034 2356 7036 2364
rect 7044 2356 7046 2364
rect 7034 2354 7046 2356
rect 7066 2804 7078 2806
rect 7066 2796 7068 2804
rect 7076 2796 7078 2804
rect 6970 1496 6972 1504
rect 6980 1496 6982 1504
rect 6344 1406 6348 1414
rect 6356 1406 6364 1414
rect 6372 1406 6380 1414
rect 6388 1406 6392 1414
rect 5946 1176 5948 1184
rect 5956 1176 5958 1184
rect 5946 1174 5958 1176
rect 5914 976 5916 984
rect 5924 976 5926 984
rect 5914 974 5926 976
rect 6344 1014 6392 1406
rect 6746 1464 6758 1466
rect 6746 1456 6748 1464
rect 6756 1456 6758 1464
rect 6746 1084 6758 1456
rect 6970 1424 6982 1496
rect 6970 1416 6972 1424
rect 6980 1416 6982 1424
rect 6970 1414 6982 1416
rect 7066 1404 7078 2796
rect 7354 2224 7366 2226
rect 7354 2216 7356 2224
rect 7364 2216 7366 2224
rect 7354 1464 7366 2216
rect 7450 1964 7462 3336
rect 7450 1956 7452 1964
rect 7460 1956 7462 1964
rect 7450 1904 7462 1956
rect 7450 1896 7452 1904
rect 7460 1896 7462 1904
rect 7450 1894 7462 1896
rect 7514 3184 7526 3186
rect 7514 3176 7516 3184
rect 7524 3176 7526 3184
rect 7514 1764 7526 3176
rect 7578 2444 7590 2446
rect 7578 2436 7580 2444
rect 7588 2436 7590 2444
rect 7578 2184 7590 2436
rect 7674 2284 7686 3936
rect 7706 3304 7718 3306
rect 7706 3296 7708 3304
rect 7716 3296 7718 3304
rect 7706 3024 7718 3296
rect 7706 3016 7708 3024
rect 7716 3016 7718 3024
rect 7706 3014 7718 3016
rect 7738 2504 7750 4056
rect 7802 3764 7814 4076
rect 7802 3756 7804 3764
rect 7812 3756 7814 3764
rect 7802 3754 7814 3756
rect 7770 3384 7782 3386
rect 7770 3376 7772 3384
rect 7780 3376 7782 3384
rect 7770 3104 7782 3376
rect 7770 3096 7772 3104
rect 7780 3096 7782 3104
rect 7770 3094 7782 3096
rect 7738 2496 7740 2504
rect 7748 2496 7750 2504
rect 7738 2494 7750 2496
rect 7770 3024 7782 3026
rect 7770 3016 7772 3024
rect 7780 3016 7782 3024
rect 7674 2276 7676 2284
rect 7684 2276 7686 2284
rect 7674 2274 7686 2276
rect 7578 2176 7580 2184
rect 7588 2176 7590 2184
rect 7578 2174 7590 2176
rect 7514 1756 7516 1764
rect 7524 1756 7526 1764
rect 7514 1754 7526 1756
rect 7706 2104 7718 2106
rect 7706 2096 7708 2104
rect 7716 2096 7718 2104
rect 7354 1456 7356 1464
rect 7364 1456 7366 1464
rect 7354 1454 7366 1456
rect 7418 1484 7430 1486
rect 7418 1476 7420 1484
rect 7428 1476 7430 1484
rect 7066 1396 7068 1404
rect 7076 1396 7078 1404
rect 7066 1394 7078 1396
rect 6746 1076 6748 1084
rect 6756 1076 6758 1084
rect 6746 1074 6758 1076
rect 6344 1006 6348 1014
rect 6356 1006 6364 1014
rect 6372 1006 6380 1014
rect 6388 1006 6392 1014
rect 6106 944 6118 946
rect 6106 936 6108 944
rect 6116 936 6118 944
rect 5466 296 5468 304
rect 5476 296 5478 304
rect 5466 294 5478 296
rect 5562 824 5574 826
rect 5562 816 5564 824
rect 5572 816 5574 824
rect 5562 164 5574 816
rect 6074 664 6086 666
rect 6074 656 6076 664
rect 6084 656 6086 664
rect 6074 524 6086 656
rect 6074 516 6076 524
rect 6084 516 6086 524
rect 6074 514 6086 516
rect 6106 284 6118 936
rect 6106 276 6108 284
rect 6116 276 6118 284
rect 6106 274 6118 276
rect 6344 614 6392 1006
rect 6344 606 6348 614
rect 6356 606 6364 614
rect 6372 606 6380 614
rect 6388 606 6392 614
rect 6344 214 6392 606
rect 7418 284 7430 1476
rect 7418 276 7420 284
rect 7428 276 7430 284
rect 7418 274 7430 276
rect 7610 844 7622 846
rect 7610 836 7612 844
rect 7620 836 7622 844
rect 7610 244 7622 836
rect 7706 844 7718 2096
rect 7770 2104 7782 3016
rect 7834 2864 7846 5096
rect 7866 3104 7878 5736
rect 8026 5724 8038 5726
rect 8026 5716 8028 5724
rect 8036 5716 8038 5724
rect 7994 5484 8006 5486
rect 7994 5476 7996 5484
rect 8004 5476 8006 5484
rect 7930 5344 7942 5346
rect 7930 5336 7932 5344
rect 7940 5336 7942 5344
rect 7898 4984 7910 4986
rect 7898 4976 7900 4984
rect 7908 4976 7910 4984
rect 7898 4864 7910 4976
rect 7898 4856 7900 4864
rect 7908 4856 7910 4864
rect 7898 4854 7910 4856
rect 7898 4164 7910 4166
rect 7898 4156 7900 4164
rect 7908 4156 7910 4164
rect 7898 3864 7910 4156
rect 7898 3856 7900 3864
rect 7908 3856 7910 3864
rect 7898 3854 7910 3856
rect 7866 3096 7868 3104
rect 7876 3096 7878 3104
rect 7866 3094 7878 3096
rect 7834 2856 7836 2864
rect 7844 2856 7846 2864
rect 7834 2854 7846 2856
rect 7930 2724 7942 5336
rect 7994 5044 8006 5476
rect 7994 5036 7996 5044
rect 8004 5036 8006 5044
rect 7994 4944 8006 5036
rect 7994 4936 7996 4944
rect 8004 4936 8006 4944
rect 7962 4764 7974 4766
rect 7962 4756 7964 4764
rect 7972 4756 7974 4764
rect 7962 3904 7974 4756
rect 7994 4444 8006 4936
rect 7994 4436 7996 4444
rect 8004 4436 8006 4444
rect 7994 4434 8006 4436
rect 7962 3896 7964 3904
rect 7972 3896 7974 3904
rect 7962 3724 7974 3896
rect 7962 3716 7964 3724
rect 7972 3716 7974 3724
rect 7962 3714 7974 3716
rect 7994 4304 8006 4306
rect 7994 4296 7996 4304
rect 8004 4296 8006 4304
rect 7994 2884 8006 4296
rect 8026 4304 8038 5716
rect 8122 5484 8134 5486
rect 8122 5476 8124 5484
rect 8132 5476 8134 5484
rect 8122 5324 8134 5476
rect 8122 5316 8124 5324
rect 8132 5316 8134 5324
rect 8122 5314 8134 5316
rect 8090 5124 8102 5126
rect 8090 5116 8092 5124
rect 8100 5116 8102 5124
rect 8058 4744 8070 4746
rect 8058 4736 8060 4744
rect 8068 4736 8070 4744
rect 8058 4664 8070 4736
rect 8058 4656 8060 4664
rect 8068 4656 8070 4664
rect 8058 4654 8070 4656
rect 8026 4296 8028 4304
rect 8036 4296 8038 4304
rect 8026 4294 8038 4296
rect 8058 4184 8070 4186
rect 8058 4176 8060 4184
rect 8068 4176 8070 4184
rect 8026 3304 8038 3306
rect 8026 3296 8028 3304
rect 8036 3296 8038 3304
rect 8026 2924 8038 3296
rect 8026 2916 8028 2924
rect 8036 2916 8038 2924
rect 8026 2914 8038 2916
rect 7994 2876 7996 2884
rect 8004 2876 8006 2884
rect 7994 2874 8006 2876
rect 7930 2716 7932 2724
rect 7940 2716 7942 2724
rect 7930 2714 7942 2716
rect 8026 2784 8038 2786
rect 8026 2776 8028 2784
rect 8036 2776 8038 2784
rect 7770 2096 7772 2104
rect 7780 2096 7782 2104
rect 7770 2094 7782 2096
rect 7802 2504 7814 2506
rect 7802 2496 7804 2504
rect 7812 2496 7814 2504
rect 7706 836 7708 844
rect 7716 836 7718 844
rect 7706 834 7718 836
rect 7802 684 7814 2496
rect 7802 676 7804 684
rect 7812 676 7814 684
rect 7802 674 7814 676
rect 7898 704 7910 706
rect 7898 696 7900 704
rect 7908 696 7910 704
rect 7898 324 7910 696
rect 8026 484 8038 2776
rect 8058 2684 8070 4176
rect 8090 3564 8102 5116
rect 8122 4924 8134 4926
rect 8122 4916 8124 4924
rect 8132 4916 8134 4924
rect 8122 4484 8134 4916
rect 8122 4476 8124 4484
rect 8132 4476 8134 4484
rect 8122 4474 8134 4476
rect 8122 4164 8134 4166
rect 8122 4156 8124 4164
rect 8132 4156 8134 4164
rect 8122 3784 8134 4156
rect 8122 3776 8124 3784
rect 8132 3776 8134 3784
rect 8122 3774 8134 3776
rect 8090 3556 8092 3564
rect 8100 3556 8102 3564
rect 8090 3554 8102 3556
rect 8058 2676 8060 2684
rect 8068 2676 8070 2684
rect 8058 2674 8070 2676
rect 8058 2604 8070 2606
rect 8058 2596 8060 2604
rect 8068 2596 8070 2604
rect 8058 744 8070 2596
rect 8058 736 8060 744
rect 8068 736 8070 744
rect 8058 734 8070 736
rect 8026 476 8028 484
rect 8036 476 8038 484
rect 8026 474 8038 476
rect 8058 524 8070 526
rect 8058 516 8060 524
rect 8068 516 8070 524
rect 7898 316 7900 324
rect 7908 316 7910 324
rect 7898 314 7910 316
rect 7962 324 7974 326
rect 7962 316 7964 324
rect 7972 316 7974 324
rect 7962 264 7974 316
rect 7962 256 7964 264
rect 7972 256 7974 264
rect 7962 254 7974 256
rect 7610 236 7612 244
rect 7620 236 7622 244
rect 7610 234 7622 236
rect 8058 244 8070 516
rect 8058 236 8060 244
rect 8068 236 8070 244
rect 8058 234 8070 236
rect 6344 206 6348 214
rect 6356 206 6364 214
rect 6372 206 6380 214
rect 6388 206 6392 214
rect 5562 156 5564 164
rect 5572 156 5574 164
rect 5562 154 5574 156
rect 5722 204 5734 206
rect 5722 196 5724 204
rect 5732 196 5734 204
rect 5722 144 5734 196
rect 5722 136 5724 144
rect 5732 136 5734 144
rect 5722 134 5734 136
rect 4808 6 4812 14
rect 4820 6 4828 14
rect 4836 6 4844 14
rect 4852 6 4856 14
rect 4808 0 4856 6
rect 6344 0 6392 206
rect 6554 154 6662 166
rect 6554 144 6566 154
rect 6554 136 6556 144
rect 6564 136 6566 144
rect 6554 134 6566 136
rect 6650 144 6662 154
rect 6650 136 6652 144
rect 6660 136 6662 144
rect 6650 134 6662 136
rect 7866 164 7878 166
rect 7866 156 7868 164
rect 7876 156 7878 164
rect 6874 124 6950 126
rect 6874 116 6876 124
rect 6884 116 6950 124
rect 6874 114 6950 116
rect 7866 124 7878 156
rect 7866 116 7868 124
rect 7876 116 7878 124
rect 7866 114 7878 116
rect 6938 104 6950 114
rect 6938 96 6940 104
rect 6948 96 6950 104
rect 6938 94 6950 96
use DFFPOSX1  DFFPOSX1_34
timestamp 1556798218
transform 1 0 8 0 -1 5810
box 0 0 192 200
use OAI21X1  OAI21X1_49
timestamp 1556798218
transform -1 0 264 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_45
timestamp 1556798218
transform -1 0 296 0 -1 5810
box 0 0 32 200
use AND2X2  AND2X2_30
timestamp 1556798218
transform -1 0 360 0 -1 5810
box 0 0 64 200
use NAND2X1  NAND2X1_65
timestamp 1556798218
transform 1 0 360 0 -1 5810
box 0 0 48 200
use INVX1  INVX1_41
timestamp 1556798218
transform -1 0 440 0 -1 5810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_39
timestamp 1556798218
transform 1 0 440 0 -1 5810
box 0 0 192 200
use INVX1  INVX1_53
timestamp 1556798218
transform 1 0 632 0 -1 5810
box 0 0 32 200
use OAI21X1  OAI21X1_57
timestamp 1556798218
transform 1 0 664 0 -1 5810
box 0 0 64 200
use CLKBUF1  CLKBUF1_24
timestamp 1556798218
transform -1 0 872 0 -1 5810
box 0 0 144 200
use NAND2X1  NAND2X1_72
timestamp 1556798218
transform 1 0 872 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_18
timestamp 1556798218
transform -1 0 1000 0 -1 5810
box 0 0 80 200
use NOR2X1  NOR2X1_32
timestamp 1556798218
transform -1 0 1048 0 -1 5810
box 0 0 48 200
use INVX1  INVX1_50
timestamp 1556798218
transform -1 0 1080 0 -1 5810
box 0 0 32 200
use NAND3X1  NAND3X1_22
timestamp 1556798218
transform -1 0 1144 0 -1 5810
box 0 0 64 200
use OAI21X1  OAI21X1_52
timestamp 1556798218
transform 1 0 1144 0 -1 5810
box 0 0 64 200
use OAI21X1  OAI21X1_53
timestamp 1556798218
transform -1 0 1272 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_49
timestamp 1556798218
transform 1 0 1272 0 -1 5810
box 0 0 32 200
use NAND3X1  NAND3X1_23
timestamp 1556798218
transform -1 0 1368 0 -1 5810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_41
timestamp 1556798218
transform 1 0 1368 0 -1 5810
box 0 0 192 200
use NAND3X1  NAND3X1_153
timestamp 1556798218
transform -1 0 1624 0 -1 5810
box 0 0 64 200
use OAI21X1  OAI21X1_450
timestamp 1556798218
transform -1 0 1688 0 -1 5810
box 0 0 64 200
use NAND2X1  NAND2X1_437
timestamp 1556798218
transform 1 0 1688 0 -1 5810
box 0 0 48 200
use FILL  FILL_28_0_0
timestamp 1556798218
transform -1 0 1752 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_0_1
timestamp 1556798218
transform -1 0 1768 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_0_2
timestamp 1556798218
transform -1 0 1784 0 -1 5810
box 0 0 16 200
use OAI21X1  OAI21X1_453
timestamp 1556798218
transform -1 0 1848 0 -1 5810
box 0 0 64 200
use CLKBUF1  CLKBUF1_12
timestamp 1556798218
transform -1 0 1992 0 -1 5810
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_298
timestamp 1556798218
transform 1 0 1992 0 -1 5810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1556798218
transform 1 0 2184 0 -1 5810
box 0 0 192 200
use OAI21X1  OAI21X1_11
timestamp 1556798218
transform -1 0 2440 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_20
timestamp 1556798218
transform -1 0 2472 0 -1 5810
box 0 0 32 200
use NAND2X1  NAND2X1_30
timestamp 1556798218
transform -1 0 2520 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_2
timestamp 1556798218
transform -1 0 2600 0 -1 5810
box 0 0 80 200
use NAND2X1  NAND2X1_31
timestamp 1556798218
transform 1 0 2600 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_3
timestamp 1556798218
transform -1 0 2728 0 -1 5810
box 0 0 80 200
use INVX1  INVX1_21
timestamp 1556798218
transform 1 0 2728 0 -1 5810
box 0 0 32 200
use OAI21X1  OAI21X1_12
timestamp 1556798218
transform 1 0 2760 0 -1 5810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1556798218
transform -1 0 3016 0 -1 5810
box 0 0 192 200
use NAND2X1  NAND2X1_33
timestamp 1556798218
transform 1 0 3016 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_5
timestamp 1556798218
transform -1 0 3144 0 -1 5810
box 0 0 80 200
use INVX1  INVX1_23
timestamp 1556798218
transform 1 0 3144 0 -1 5810
box 0 0 32 200
use OAI21X1  OAI21X1_14
timestamp 1556798218
transform 1 0 3176 0 -1 5810
box 0 0 64 200
use FILL  FILL_28_1_0
timestamp 1556798218
transform -1 0 3256 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_1_1
timestamp 1556798218
transform -1 0 3272 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_1_2
timestamp 1556798218
transform -1 0 3288 0 -1 5810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1556798218
transform -1 0 3480 0 -1 5810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1556798218
transform 1 0 3480 0 -1 5810
box 0 0 192 200
use INVX1  INVX1_24
timestamp 1556798218
transform 1 0 3672 0 -1 5810
box 0 0 32 200
use OAI21X1  OAI21X1_15
timestamp 1556798218
transform 1 0 3704 0 -1 5810
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1556798218
transform -1 0 3816 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_6
timestamp 1556798218
transform -1 0 3896 0 -1 5810
box 0 0 80 200
use BUFX2  BUFX2_135
timestamp 1556798218
transform 1 0 3896 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_1
timestamp 1556798218
transform 1 0 3944 0 -1 5810
box 0 0 80 200
use NAND2X1  NAND2X1_29
timestamp 1556798218
transform 1 0 4024 0 -1 5810
box 0 0 48 200
use OAI21X1  OAI21X1_10
timestamp 1556798218
transform -1 0 4136 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_18
timestamp 1556798218
transform -1 0 4168 0 -1 5810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1556798218
transform -1 0 4360 0 -1 5810
box 0 0 192 200
use INVX1  INVX1_15
timestamp 1556798218
transform -1 0 4392 0 -1 5810
box 0 0 32 200
use XNOR2X1  XNOR2X1_69
timestamp 1556798218
transform 1 0 4392 0 -1 5810
box 0 0 112 200
use AOI21X1  AOI21X1_74
timestamp 1556798218
transform 1 0 4504 0 -1 5810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_304
timestamp 1556798218
transform 1 0 4568 0 -1 5810
box 0 0 192 200
use INVX1  INVX1_513
timestamp 1556798218
transform -1 0 4792 0 -1 5810
box 0 0 32 200
use FILL  FILL_28_2_0
timestamp 1556798218
transform -1 0 4808 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_2_1
timestamp 1556798218
transform -1 0 4824 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_2_2
timestamp 1556798218
transform -1 0 4840 0 -1 5810
box 0 0 16 200
use CLKBUF1  CLKBUF1_21
timestamp 1556798218
transform -1 0 4984 0 -1 5810
box 0 0 144 200
use AND2X2  AND2X2_120
timestamp 1556798218
transform 1 0 4984 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_528
timestamp 1556798218
transform 1 0 5048 0 -1 5810
box 0 0 32 200
use NAND2X1  NAND2X1_451
timestamp 1556798218
transform 1 0 5080 0 -1 5810
box 0 0 48 200
use OAI21X1  OAI21X1_470
timestamp 1556798218
transform 1 0 5128 0 -1 5810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_310
timestamp 1556798218
transform 1 0 5192 0 -1 5810
box 0 0 192 200
use NAND2X1  NAND2X1_455
timestamp 1556798218
transform 1 0 5384 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_155
timestamp 1556798218
transform 1 0 5432 0 -1 5810
box 0 0 80 200
use OAI21X1  OAI21X1_469
timestamp 1556798218
transform -1 0 5576 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_527
timestamp 1556798218
transform 1 0 5576 0 -1 5810
box 0 0 32 200
use NOR2X1  NOR2X1_204
timestamp 1556798218
transform 1 0 5608 0 -1 5810
box 0 0 48 200
use INVX1  INVX1_526
timestamp 1556798218
transform -1 0 5688 0 -1 5810
box 0 0 32 200
use AOI21X1  AOI21X1_76
timestamp 1556798218
transform 1 0 5688 0 -1 5810
box 0 0 64 200
use NAND3X1  NAND3X1_158
timestamp 1556798218
transform -1 0 5816 0 -1 5810
box 0 0 64 200
use NAND2X1  NAND2X1_453
timestamp 1556798218
transform -1 0 5864 0 -1 5810
box 0 0 48 200
use AOI22X1  AOI22X1_154
timestamp 1556798218
transform -1 0 5944 0 -1 5810
box 0 0 80 200
use XNOR2X1  XNOR2X1_71
timestamp 1556798218
transform -1 0 6056 0 -1 5810
box 0 0 112 200
use OAI21X1  OAI21X1_472
timestamp 1556798218
transform -1 0 6120 0 -1 5810
box 0 0 64 200
use INVX1  INVX1_529
timestamp 1556798218
transform -1 0 6152 0 -1 5810
box 0 0 32 200
use BUFX2  BUFX2_4
timestamp 1556798218
transform 1 0 6152 0 -1 5810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_311
timestamp 1556798218
transform -1 0 6392 0 -1 5810
box 0 0 192 200
use FILL  FILL_28_3_0
timestamp 1556798218
transform -1 0 6408 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_3_1
timestamp 1556798218
transform -1 0 6424 0 -1 5810
box 0 0 16 200
use FILL  FILL_28_3_2
timestamp 1556798218
transform -1 0 6440 0 -1 5810
box 0 0 16 200
use CLKBUF1  CLKBUF1_51
timestamp 1556798218
transform -1 0 6584 0 -1 5810
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_50
timestamp 1556798218
transform -1 0 6776 0 -1 5810
box 0 0 192 200
use CLKBUF1  CLKBUF1_22
timestamp 1556798218
transform 1 0 6776 0 -1 5810
box 0 0 144 200
use NAND3X1  NAND3X1_163
timestamp 1556798218
transform -1 0 6984 0 -1 5810
box 0 0 64 200
use OAI21X1  OAI21X1_480
timestamp 1556798218
transform -1 0 7048 0 -1 5810
box 0 0 64 200
use NAND2X1  NAND2X1_462
timestamp 1556798218
transform 1 0 7048 0 -1 5810
box 0 0 48 200
use OAI21X1  OAI21X1_483
timestamp 1556798218
transform -1 0 7160 0 -1 5810
box 0 0 64 200
use AOI21X1  AOI21X1_78
timestamp 1556798218
transform -1 0 7224 0 -1 5810
box 0 0 64 200
use XNOR2X1  XNOR2X1_73
timestamp 1556798218
transform -1 0 7336 0 -1 5810
box 0 0 112 200
use XNOR2X1  XNOR2X1_34
timestamp 1556798218
transform 1 0 7336 0 -1 5810
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_168
timestamp 1556798218
transform -1 0 7640 0 -1 5810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_176
timestamp 1556798218
transform 1 0 7640 0 -1 5810
box 0 0 192 200
use CLKBUF1  CLKBUF1_28
timestamp 1556798218
transform 1 0 7832 0 -1 5810
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1556798218
transform 1 0 7976 0 -1 5810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_37
timestamp 1556798218
transform 1 0 8 0 1 5410
box 0 0 192 200
use AOI22X1  AOI22X1_17
timestamp 1556798218
transform -1 0 280 0 1 5410
box 0 0 80 200
use NOR2X1  NOR2X1_30
timestamp 1556798218
transform -1 0 328 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_48
timestamp 1556798218
transform -1 0 392 0 1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_69
timestamp 1556798218
transform -1 0 440 0 1 5410
box 0 0 48 200
use INVX1  INVX1_44
timestamp 1556798218
transform 1 0 440 0 1 5410
box 0 0 32 200
use NAND3X1  NAND3X1_21
timestamp 1556798218
transform 1 0 472 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_20
timestamp 1556798218
transform 1 0 536 0 1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_29
timestamp 1556798218
transform 1 0 600 0 1 5410
box 0 0 48 200
use INVX1  INVX1_40
timestamp 1556798218
transform -1 0 680 0 1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_36
timestamp 1556798218
transform -1 0 872 0 1 5410
box 0 0 192 200
use AND2X2  AND2X2_29
timestamp 1556798218
transform 1 0 872 0 1 5410
box 0 0 64 200
use INVX1  INVX1_51
timestamp 1556798218
transform 1 0 936 0 1 5410
box 0 0 32 200
use AOI22X1  AOI22X1_19
timestamp 1556798218
transform 1 0 968 0 1 5410
box 0 0 80 200
use NAND2X1  NAND2X1_74
timestamp 1556798218
transform 1 0 1048 0 1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_73
timestamp 1556798218
transform -1 0 1144 0 1 5410
box 0 0 48 200
use INVX1  INVX1_48
timestamp 1556798218
transform -1 0 1176 0 1 5410
box 0 0 32 200
use AOI21X1  AOI21X1_8
timestamp 1556798218
transform 1 0 1176 0 1 5410
box 0 0 64 200
use AND2X2  AND2X2_31
timestamp 1556798218
transform -1 0 1304 0 1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_71
timestamp 1556798218
transform 1 0 1304 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_54
timestamp 1556798218
transform 1 0 1352 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_56
timestamp 1556798218
transform 1 0 1416 0 1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_31
timestamp 1556798218
transform 1 0 1480 0 1 5410
box 0 0 48 200
use INVX1  INVX1_47
timestamp 1556798218
transform -1 0 1560 0 1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_301
timestamp 1556798218
transform 1 0 1560 0 1 5410
box 0 0 192 200
use FILL  FILL_27_0_0
timestamp 1556798218
transform -1 0 1768 0 1 5410
box 0 0 16 200
use FILL  FILL_27_0_1
timestamp 1556798218
transform -1 0 1784 0 1 5410
box 0 0 16 200
use FILL  FILL_27_0_2
timestamp 1556798218
transform -1 0 1800 0 1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_73
timestamp 1556798218
transform -1 0 1864 0 1 5410
box 0 0 64 200
use INVX1  INVX1_504
timestamp 1556798218
transform 1 0 1864 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_449
timestamp 1556798218
transform -1 0 1960 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_152
timestamp 1556798218
transform 1 0 1960 0 1 5410
box 0 0 64 200
use INVX1  INVX1_506
timestamp 1556798218
transform 1 0 2024 0 1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_438
timestamp 1556798218
transform -1 0 2104 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_451
timestamp 1556798218
transform 1 0 2104 0 1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_436
timestamp 1556798218
transform 1 0 2168 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_452
timestamp 1556798218
transform -1 0 2280 0 1 5410
box 0 0 64 200
use INVX1  INVX1_507
timestamp 1556798218
transform -1 0 2312 0 1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_197
timestamp 1556798218
transform 1 0 2312 0 1 5410
box 0 0 48 200
use INVX1  INVX1_502
timestamp 1556798218
transform -1 0 2392 0 1 5410
box 0 0 32 200
use BUFX2  BUFX2_29
timestamp 1556798218
transform -1 0 2440 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_7
timestamp 1556798218
transform -1 0 2488 0 1 5410
box 0 0 48 200
use CLKBUF1  CLKBUF1_34
timestamp 1556798218
transform 1 0 2488 0 1 5410
box 0 0 144 200
use NAND2X1  NAND2X1_32
timestamp 1556798218
transform -1 0 2680 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_13
timestamp 1556798218
transform -1 0 2744 0 1 5410
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1556798218
transform -1 0 2776 0 1 5410
box 0 0 32 200
use AOI22X1  AOI22X1_4
timestamp 1556798218
transform 1 0 2776 0 1 5410
box 0 0 80 200
use NAND2X1  NAND2X1_38
timestamp 1556798218
transform -1 0 2904 0 1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_39
timestamp 1556798218
transform -1 0 2952 0 1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1556798218
transform 1 0 2952 0 1 5410
box 0 0 192 200
use NAND2X1  NAND2X1_41
timestamp 1556798218
transform -1 0 3192 0 1 5410
box 0 0 48 200
use FILL  FILL_27_1_0
timestamp 1556798218
transform 1 0 3192 0 1 5410
box 0 0 16 200
use FILL  FILL_27_1_1
timestamp 1556798218
transform 1 0 3208 0 1 5410
box 0 0 16 200
use FILL  FILL_27_1_2
timestamp 1556798218
transform 1 0 3224 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1556798218
transform 1 0 3240 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_16
timestamp 1556798218
transform -1 0 3496 0 1 5410
box 0 0 64 200
use INVX1  INVX1_25
timestamp 1556798218
transform -1 0 3528 0 1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_35
timestamp 1556798218
transform -1 0 3576 0 1 5410
box 0 0 48 200
use AOI22X1  AOI22X1_7
timestamp 1556798218
transform 1 0 3576 0 1 5410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1556798218
transform 1 0 3656 0 1 5410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1556798218
transform -1 0 4040 0 1 5410
box 0 0 192 200
use NAND2X1  NAND2X1_37
timestamp 1556798218
transform -1 0 4088 0 1 5410
box 0 0 48 200
use NOR2X1  NOR2X1_19
timestamp 1556798218
transform 1 0 4088 0 1 5410
box 0 0 48 200
use INVX1  INVX1_19
timestamp 1556798218
transform -1 0 4168 0 1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_17
timestamp 1556798218
transform -1 0 4216 0 1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_36
timestamp 1556798218
transform -1 0 4264 0 1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_28
timestamp 1556798218
transform 1 0 4264 0 1 5410
box 0 0 48 200
use INVX1  INVX1_17
timestamp 1556798218
transform -1 0 4344 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_8
timestamp 1556798218
transform -1 0 4408 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1556798218
transform -1 0 4472 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_19
timestamp 1556798218
transform 1 0 4472 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_14
timestamp 1556798218
transform 1 0 4536 0 1 5410
box 0 0 64 200
use CLKBUF1  CLKBUF1_18
timestamp 1556798218
transform -1 0 4744 0 1 5410
box 0 0 144 200
use INVX1  INVX1_511
timestamp 1556798218
transform 1 0 4744 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_459
timestamp 1556798218
transform -1 0 4840 0 1 5410
box 0 0 64 200
use FILL  FILL_27_2_0
timestamp 1556798218
transform 1 0 4840 0 1 5410
box 0 0 16 200
use FILL  FILL_27_2_1
timestamp 1556798218
transform 1 0 4856 0 1 5410
box 0 0 16 200
use FILL  FILL_27_2_2
timestamp 1556798218
transform 1 0 4872 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_442
timestamp 1556798218
transform 1 0 4888 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_455
timestamp 1556798218
transform -1 0 5000 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_154
timestamp 1556798218
transform 1 0 5000 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_456
timestamp 1556798218
transform -1 0 5128 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_155
timestamp 1556798218
transform 1 0 5128 0 1 5410
box 0 0 64 200
use INVX1  INVX1_512
timestamp 1556798218
transform -1 0 5224 0 1 5410
box 0 0 32 200
use BUFX2  BUFX2_63
timestamp 1556798218
transform -1 0 5272 0 1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_305
timestamp 1556798218
transform -1 0 5464 0 1 5410
box 0 0 192 200
use NOR2X1  NOR2X1_192
timestamp 1556798218
transform -1 0 5512 0 1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_454
timestamp 1556798218
transform -1 0 5560 0 1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_312
timestamp 1556798218
transform 1 0 5560 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_468
timestamp 1556798218
transform 1 0 5752 0 1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_159
timestamp 1556798218
transform -1 0 5880 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_467
timestamp 1556798218
transform 1 0 5880 0 1 5410
box 0 0 64 200
use INVX1  INVX1_525
timestamp 1556798218
transform 1 0 5944 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_471
timestamp 1556798218
transform 1 0 5976 0 1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_452
timestamp 1556798218
transform 1 0 6040 0 1 5410
box 0 0 48 200
use INVX1  INVX1_524
timestamp 1556798218
transform -1 0 6120 0 1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_203
timestamp 1556798218
transform 1 0 6120 0 1 5410
box 0 0 48 200
use INVX1  INVX1_523
timestamp 1556798218
transform -1 0 6200 0 1 5410
box 0 0 32 200
use AND2X2  AND2X2_13
timestamp 1556798218
transform 1 0 6200 0 1 5410
box 0 0 64 200
use AOI21X1  AOI21X1_11
timestamp 1556798218
transform -1 0 6328 0 1 5410
box 0 0 64 200
use FILL  FILL_27_3_0
timestamp 1556798218
transform -1 0 6344 0 1 5410
box 0 0 16 200
use FILL  FILL_27_3_1
timestamp 1556798218
transform -1 0 6360 0 1 5410
box 0 0 16 200
use FILL  FILL_27_3_2
timestamp 1556798218
transform -1 0 6376 0 1 5410
box 0 0 16 200
use XNOR2X1  XNOR2X1_6
timestamp 1556798218
transform -1 0 6488 0 1 5410
box 0 0 112 200
use AND2X2  AND2X2_34
timestamp 1556798218
transform 1 0 6488 0 1 5410
box 0 0 64 200
use AOI22X1  AOI22X1_25
timestamp 1556798218
transform 1 0 6552 0 1 5410
box 0 0 80 200
use OAI21X1  OAI21X1_73
timestamp 1556798218
transform 1 0 6632 0 1 5410
box 0 0 64 200
use INVX1  INVX1_73
timestamp 1556798218
transform 1 0 6696 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_74
timestamp 1556798218
transform 1 0 6728 0 1 5410
box 0 0 64 200
use BUFX2  BUFX2_66
timestamp 1556798218
transform -1 0 6840 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_64
timestamp 1556798218
transform 1 0 6840 0 1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_321
timestamp 1556798218
transform 1 0 6888 0 1 5410
box 0 0 192 200
use INVX1  INVX1_538
timestamp 1556798218
transform 1 0 7080 0 1 5410
box 0 0 32 200
use NAND3X1  NAND3X1_162
timestamp 1556798218
transform 1 0 7112 0 1 5410
box 0 0 64 200
use INVX1  INVX1_537
timestamp 1556798218
transform 1 0 7176 0 1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_207
timestamp 1556798218
transform -1 0 7256 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_479
timestamp 1556798218
transform 1 0 7256 0 1 5410
box 0 0 64 200
use INVX1  INVX1_539
timestamp 1556798218
transform -1 0 7352 0 1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_320
timestamp 1556798218
transform -1 0 7544 0 1 5410
box 0 0 192 200
use INVX1  INVX1_285
timestamp 1556798218
transform 1 0 7544 0 1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_104
timestamp 1556798218
transform -1 0 7624 0 1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_177
timestamp 1556798218
transform -1 0 7816 0 1 5410
box 0 0 192 200
use INVX1  INVX1_286
timestamp 1556798218
transform 1 0 7816 0 1 5410
box 0 0 32 200
use NAND3X1  NAND3X1_91
timestamp 1556798218
transform 1 0 7848 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_263
timestamp 1556798218
transform -1 0 7976 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_262
timestamp 1556798218
transform 1 0 7976 0 1 5410
box 0 0 64 200
use INVX1  INVX1_287
timestamp 1556798218
transform 1 0 8040 0 1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_266
timestamp 1556798218
transform -1 0 8136 0 1 5410
box 0 0 64 200
use FILL  FILL_28_1
timestamp 1556798218
transform 1 0 8136 0 1 5410
box 0 0 16 200
use FILL  FILL_28_2
timestamp 1556798218
transform 1 0 8152 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_35
timestamp 1556798218
transform -1 0 200 0 -1 5410
box 0 0 192 200
use INVX1  INVX1_46
timestamp 1556798218
transform 1 0 200 0 -1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_51
timestamp 1556798218
transform -1 0 296 0 -1 5410
box 0 0 64 200
use AOI22X1  AOI22X1_16
timestamp 1556798218
transform -1 0 376 0 -1 5410
box 0 0 80 200
use NAND2X1  NAND2X1_67
timestamp 1556798218
transform -1 0 424 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_68
timestamp 1556798218
transform -1 0 472 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_47
timestamp 1556798218
transform 1 0 472 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_46
timestamp 1556798218
transform 1 0 536 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_42
timestamp 1556798218
transform -1 0 632 0 -1 5410
box 0 0 32 200
use INVX1  INVX1_43
timestamp 1556798218
transform -1 0 664 0 -1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_66
timestamp 1556798218
transform -1 0 712 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_50
timestamp 1556798218
transform 1 0 712 0 -1 5410
box 0 0 64 200
use AOI21X1  AOI21X1_7
timestamp 1556798218
transform -1 0 840 0 -1 5410
box 0 0 64 200
use XNOR2X1  XNOR2X1_2
timestamp 1556798218
transform -1 0 952 0 -1 5410
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_40
timestamp 1556798218
transform 1 0 952 0 -1 5410
box 0 0 192 200
use XNOR2X1  XNOR2X1_3
timestamp 1556798218
transform 1 0 1144 0 -1 5410
box 0 0 112 200
use NAND2X1  NAND2X1_70
timestamp 1556798218
transform -1 0 1304 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_52
timestamp 1556798218
transform 1 0 1304 0 -1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_55
timestamp 1556798218
transform 1 0 1336 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_38
timestamp 1556798218
transform -1 0 1592 0 -1 5410
box 0 0 192 200
use NOR2X1  NOR2X1_44
timestamp 1556798218
transform 1 0 1592 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_89
timestamp 1556798218
transform 1 0 1640 0 -1 5410
box 0 0 32 200
use INVX1  INVX1_503
timestamp 1556798218
transform -1 0 1704 0 -1 5410
box 0 0 32 200
use BUFX2  BUFX2_23
timestamp 1556798218
transform 1 0 1704 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_0_0
timestamp 1556798218
transform -1 0 1768 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_0_1
timestamp 1556798218
transform -1 0 1784 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_0_2
timestamp 1556798218
transform -1 0 1800 0 -1 5410
box 0 0 16 200
use XNOR2X1  XNOR2X1_68
timestamp 1556798218
transform -1 0 1912 0 -1 5410
box 0 0 112 200
use BUFX2  BUFX2_25
timestamp 1556798218
transform 1 0 1912 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_505
timestamp 1556798218
transform 1 0 1960 0 -1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_198
timestamp 1556798218
transform 1 0 1992 0 -1 5410
box 0 0 48 200
use AOI22X1  AOI22X1_148
timestamp 1556798218
transform -1 0 2120 0 -1 5410
box 0 0 80 200
use AND2X2  AND2X2_117
timestamp 1556798218
transform 1 0 2120 0 -1 5410
box 0 0 64 200
use AOI22X1  AOI22X1_149
timestamp 1556798218
transform -1 0 2264 0 -1 5410
box 0 0 80 200
use NAND2X1  NAND2X1_439
timestamp 1556798218
transform 1 0 2264 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_440
timestamp 1556798218
transform -1 0 2360 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_454
timestamp 1556798218
transform -1 0 2424 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_299
timestamp 1556798218
transform 1 0 2424 0 -1 5410
box 0 0 192 200
use INVX1  INVX1_508
timestamp 1556798218
transform -1 0 2648 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1556798218
transform 1 0 2648 0 -1 5410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1556798218
transform 1 0 2840 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_20
timestamp 1556798218
transform -1 0 3096 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_21
timestamp 1556798218
transform -1 0 3160 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_23
timestamp 1556798218
transform 1 0 3160 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_9
timestamp 1556798218
transform 1 0 3224 0 -1 5410
box 0 0 32 200
use FILL  FILL_26_1_0
timestamp 1556798218
transform 1 0 3256 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_1_1
timestamp 1556798218
transform 1 0 3272 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_1_2
timestamp 1556798218
transform 1 0 3288 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1556798218
transform 1 0 3304 0 -1 5410
box 0 0 192 200
use NAND2X1  NAND2X1_40
timestamp 1556798218
transform -1 0 3544 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_22
timestamp 1556798218
transform 1 0 3544 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_43
timestamp 1556798218
transform -1 0 3656 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_25
timestamp 1556798218
transform 1 0 3656 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1556798218
transform 1 0 3720 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_18
timestamp 1556798218
transform -1 0 3976 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_18
timestamp 1556798218
transform -1 0 4024 0 -1 5410
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1556798218
transform -1 0 4088 0 -1 5410
box 0 0 64 200
use AOI21X1  AOI21X1_1
timestamp 1556798218
transform 1 0 4088 0 -1 5410
box 0 0 64 200
use AND2X2  AND2X2_23
timestamp 1556798218
transform -1 0 4216 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_17
timestamp 1556798218
transform 1 0 4216 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_16
timestamp 1556798218
transform 1 0 4280 0 -1 5410
box 0 0 32 200
use OR2X2  OR2X2_1
timestamp 1556798218
transform 1 0 4312 0 -1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_13
timestamp 1556798218
transform 1 0 4376 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1556798218
transform 1 0 4440 0 -1 5410
box 0 0 192 200
use CLKBUF1  CLKBUF1_5
timestamp 1556798218
transform -1 0 4776 0 -1 5410
box 0 0 144 200
use NOR2X1  NOR2X1_199
timestamp 1556798218
transform -1 0 4824 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_2_0
timestamp 1556798218
transform -1 0 4840 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_2_1
timestamp 1556798218
transform -1 0 4856 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_2_2
timestamp 1556798218
transform -1 0 4872 0 -1 5410
box 0 0 16 200
use OAI21X1  OAI21X1_457
timestamp 1556798218
transform -1 0 4936 0 -1 5410
box 0 0 64 200
use BUFX2  BUFX2_89
timestamp 1556798218
transform 1 0 4936 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_510
timestamp 1556798218
transform 1 0 4984 0 -1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_443
timestamp 1556798218
transform 1 0 5016 0 -1 5410
box 0 0 48 200
use AOI22X1  AOI22X1_150
timestamp 1556798218
transform -1 0 5144 0 -1 5410
box 0 0 80 200
use NOR2X1  NOR2X1_200
timestamp 1556798218
transform -1 0 5192 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_444
timestamp 1556798218
transform -1 0 5240 0 -1 5410
box 0 0 48 200
use BUFX2  BUFX2_61
timestamp 1556798218
transform -1 0 5288 0 -1 5410
box 0 0 48 200
use NOR2X1  NOR2X1_195
timestamp 1556798218
transform 1 0 5288 0 -1 5410
box 0 0 48 200
use NOR2X1  NOR2X1_196
timestamp 1556798218
transform 1 0 5336 0 -1 5410
box 0 0 48 200
use AND2X2  AND2X2_116
timestamp 1556798218
transform -1 0 5448 0 -1 5410
box 0 0 64 200
use AND2X2  AND2X2_114
timestamp 1556798218
transform -1 0 5512 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_191
timestamp 1556798218
transform -1 0 5560 0 -1 5410
box 0 0 48 200
use CLKBUF1  CLKBUF1_26
timestamp 1556798218
transform 1 0 5560 0 -1 5410
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_313
timestamp 1556798218
transform -1 0 5896 0 -1 5410
box 0 0 192 200
use INVX1  INVX1_68
timestamp 1556798218
transform 1 0 5896 0 -1 5410
box 0 0 32 200
use NOR2X1  NOR2X1_37
timestamp 1556798218
transform -1 0 5976 0 -1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_52
timestamp 1556798218
transform 1 0 5976 0 -1 5410
box 0 0 192 200
use NAND3X1  NAND3X1_29
timestamp 1556798218
transform -1 0 6232 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_75
timestamp 1556798218
transform -1 0 6296 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_70
timestamp 1556798218
transform -1 0 6328 0 -1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_88
timestamp 1556798218
transform -1 0 6376 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_3_0
timestamp 1556798218
transform 1 0 6376 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_3_1
timestamp 1556798218
transform 1 0 6392 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_3_2
timestamp 1556798218
transform 1 0 6408 0 -1 5410
box 0 0 16 200
use NAND3X1  NAND3X1_28
timestamp 1556798218
transform 1 0 6424 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_90
timestamp 1556798218
transform -1 0 6536 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_91
timestamp 1556798218
transform -1 0 6584 0 -1 5410
box 0 0 48 200
use NOR2X1  NOR2X1_38
timestamp 1556798218
transform 1 0 6584 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_69
timestamp 1556798218
transform -1 0 6664 0 -1 5410
box 0 0 32 200
use NAND2X1  NAND2X1_87
timestamp 1556798218
transform 1 0 6664 0 -1 5410
box 0 0 48 200
use AND2X2  AND2X2_122
timestamp 1556798218
transform 1 0 6712 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_542
timestamp 1556798218
transform 1 0 6776 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_318
timestamp 1556798218
transform 1 0 6808 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_482
timestamp 1556798218
transform 1 0 7000 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_461
timestamp 1556798218
transform 1 0 7064 0 -1 5410
box 0 0 48 200
use AOI22X1  AOI22X1_159
timestamp 1556798218
transform 1 0 7112 0 -1 5410
box 0 0 80 200
use OAI21X1  OAI21X1_481
timestamp 1556798218
transform -1 0 7256 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_463
timestamp 1556798218
transform 1 0 7256 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_541
timestamp 1556798218
transform -1 0 7336 0 -1 5410
box 0 0 32 200
use AOI22X1  AOI22X1_158
timestamp 1556798218
transform 1 0 7336 0 -1 5410
box 0 0 80 200
use NOR2X1  NOR2X1_208
timestamp 1556798218
transform 1 0 7416 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_540
timestamp 1556798218
transform -1 0 7496 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_174
timestamp 1556798218
transform 1 0 7496 0 -1 5410
box 0 0 192 200
use AOI22X1  AOI22X1_86
timestamp 1556798218
transform 1 0 7688 0 -1 5410
box 0 0 80 200
use NAND2X1  NAND2X1_264
timestamp 1556798218
transform 1 0 7768 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_264
timestamp 1556798218
transform -1 0 7880 0 -1 5410
box 0 0 64 200
use NAND3X1  NAND3X1_90
timestamp 1556798218
transform 1 0 7880 0 -1 5410
box 0 0 64 200
use INVX1  INVX1_288
timestamp 1556798218
transform -1 0 7976 0 -1 5410
box 0 0 32 200
use AOI21X1  AOI21X1_42
timestamp 1556798218
transform 1 0 7976 0 -1 5410
box 0 0 64 200
use XNOR2X1  XNOR2X1_37
timestamp 1556798218
transform -1 0 8152 0 -1 5410
box 0 0 112 200
use FILL  FILL_27_1
timestamp 1556798218
transform -1 0 8168 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_88
timestamp 1556798218
transform 1 0 8 0 1 5010
box 0 0 192 200
use AOI21X1  AOI21X1_20
timestamp 1556798218
transform -1 0 264 0 1 5010
box 0 0 64 200
use XNOR2X1  XNOR2X1_15
timestamp 1556798218
transform -1 0 376 0 1 5010
box 0 0 112 200
use NOR2X1  NOR2X1_57
timestamp 1556798218
transform 1 0 376 0 1 5010
box 0 0 48 200
use INVX1  INVX1_131
timestamp 1556798218
transform -1 0 456 0 1 5010
box 0 0 32 200
use BUFX2  BUFX2_24
timestamp 1556798218
transform -1 0 504 0 1 5010
box 0 0 48 200
use INVX1  INVX1_135
timestamp 1556798218
transform -1 0 536 0 1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_1
timestamp 1556798218
transform -1 0 584 0 1 5010
box 0 0 48 200
use NOR2X1  NOR2X1_1
timestamp 1556798218
transform 1 0 584 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_2
timestamp 1556798218
transform 1 0 632 0 1 5010
box 0 0 48 200
use CLKBUF1  CLKBUF1_2
timestamp 1556798218
transform -1 0 824 0 1 5010
box 0 0 144 200
use BUFX2  BUFX2_50
timestamp 1556798218
transform -1 0 872 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_56
timestamp 1556798218
transform 1 0 872 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_64
timestamp 1556798218
transform 1 0 920 0 1 5010
box 0 0 192 200
use AOI21X1  AOI21X1_14
timestamp 1556798218
transform 1 0 1112 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_93
timestamp 1556798218
transform -1 0 1240 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_106
timestamp 1556798218
transform 1 0 1240 0 1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_34
timestamp 1556798218
transform -1 0 1352 0 1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_35
timestamp 1556798218
transform 1 0 1352 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_65
timestamp 1556798218
transform 1 0 1416 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_300
timestamp 1556798218
transform 1 0 1608 0 1 5010
box 0 0 192 200
use FILL  FILL_25_0_0
timestamp 1556798218
transform 1 0 1800 0 1 5010
box 0 0 16 200
use FILL  FILL_25_0_1
timestamp 1556798218
transform 1 0 1816 0 1 5010
box 0 0 16 200
use FILL  FILL_25_0_2
timestamp 1556798218
transform 1 0 1832 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_136
timestamp 1556798218
transform 1 0 1848 0 1 5010
box 0 0 192 200
use INVX1  INVX1_215
timestamp 1556798218
transform 1 0 2040 0 1 5010
box 0 0 32 200
use NOR2X1  NOR2X1_83
timestamp 1556798218
transform -1 0 2120 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_204
timestamp 1556798218
transform -1 0 2184 0 1 5010
box 0 0 64 200
use AOI21X1  AOI21X1_32
timestamp 1556798218
transform -1 0 2248 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_207
timestamp 1556798218
transform -1 0 2296 0 1 5010
box 0 0 48 200
use XNOR2X1  XNOR2X1_27
timestamp 1556798218
transform 1 0 2296 0 1 5010
box 0 0 112 200
use INVX1  INVX1_219
timestamp 1556798218
transform -1 0 2440 0 1 5010
box 0 0 32 200
use INVX1  INVX1_216
timestamp 1556798218
transform 1 0 2440 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_202
timestamp 1556798218
transform 1 0 2472 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_206
timestamp 1556798218
transform 1 0 2536 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_203
timestamp 1556798218
transform -1 0 2648 0 1 5010
box 0 0 64 200
use INVX1  INVX1_220
timestamp 1556798218
transform -1 0 2680 0 1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_134
timestamp 1556798218
transform 1 0 2680 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_210
timestamp 1556798218
transform 1 0 2872 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_209
timestamp 1556798218
transform -1 0 2968 0 1 5010
box 0 0 48 200
use AND2X2  AND2X2_57
timestamp 1556798218
transform -1 0 3032 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_130
timestamp 1556798218
transform 1 0 3032 0 1 5010
box 0 0 192 200
use INVX1  INVX1_213
timestamp 1556798218
transform 1 0 3224 0 1 5010
box 0 0 32 200
use FILL  FILL_25_1_0
timestamp 1556798218
transform 1 0 3256 0 1 5010
box 0 0 16 200
use FILL  FILL_25_1_1
timestamp 1556798218
transform 1 0 3272 0 1 5010
box 0 0 16 200
use FILL  FILL_25_1_2
timestamp 1556798218
transform 1 0 3288 0 1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_197
timestamp 1556798218
transform 1 0 3304 0 1 5010
box 0 0 64 200
use AND2X2  AND2X2_58
timestamp 1556798218
transform 1 0 3368 0 1 5010
box 0 0 64 200
use AOI22X1  AOI22X1_65
timestamp 1556798218
transform 1 0 3432 0 1 5010
box 0 0 80 200
use OAI21X1  OAI21X1_196
timestamp 1556798218
transform -1 0 3576 0 1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_82
timestamp 1556798218
transform -1 0 3624 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_203
timestamp 1556798218
transform -1 0 3672 0 1 5010
box 0 0 48 200
use AOI22X1  AOI22X1_64
timestamp 1556798218
transform 1 0 3672 0 1 5010
box 0 0 80 200
use OAI21X1  OAI21X1_199
timestamp 1556798218
transform -1 0 3816 0 1 5010
box 0 0 64 200
use INVX1  INVX1_214
timestamp 1556798218
transform -1 0 3848 0 1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_42
timestamp 1556798218
transform -1 0 3896 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1556798218
transform 1 0 3896 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_131
timestamp 1556798218
transform 1 0 3960 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1556798218
transform 1 0 4152 0 1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_16
timestamp 1556798218
transform 1 0 4344 0 1 5010
box 0 0 48 200
use INVX1  INVX1_14
timestamp 1556798218
transform -1 0 4424 0 1 5010
box 0 0 32 200
use INVX1  INVX1_509
timestamp 1556798218
transform 1 0 4424 0 1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_302
timestamp 1556798218
transform 1 0 4456 0 1 5010
box 0 0 192 200
use INVX1  INVX1_514
timestamp 1556798218
transform 1 0 4648 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_458
timestamp 1556798218
transform 1 0 4680 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_441
timestamp 1556798218
transform -1 0 4792 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_433
timestamp 1556798218
transform 1 0 4792 0 1 5010
box 0 0 48 200
use FILL  FILL_25_2_0
timestamp 1556798218
transform -1 0 4856 0 1 5010
box 0 0 16 200
use FILL  FILL_25_2_1
timestamp 1556798218
transform -1 0 4872 0 1 5010
box 0 0 16 200
use FILL  FILL_25_2_2
timestamp 1556798218
transform -1 0 4888 0 1 5010
box 0 0 16 200
use AOI22X1  AOI22X1_151
timestamp 1556798218
transform -1 0 4968 0 1 5010
box 0 0 80 200
use NAND2X1  NAND2X1_445
timestamp 1556798218
transform 1 0 4968 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_460
timestamp 1556798218
transform -1 0 5080 0 1 5010
box 0 0 64 200
use INVX1  INVX1_515
timestamp 1556798218
transform -1 0 5112 0 1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_303
timestamp 1556798218
transform 1 0 5112 0 1 5010
box 0 0 192 200
use INVX1  INVX1_61
timestamp 1556798218
transform 1 0 5304 0 1 5010
box 0 0 32 200
use NOR2X1  NOR2X1_35
timestamp 1556798218
transform -1 0 5384 0 1 5010
box 0 0 48 200
use NOR2X1  NOR2X1_193
timestamp 1556798218
transform -1 0 5432 0 1 5010
box 0 0 48 200
use AND2X2  AND2X2_115
timestamp 1556798218
transform 1 0 5432 0 1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_194
timestamp 1556798218
transform -1 0 5544 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_47
timestamp 1556798218
transform 1 0 5544 0 1 5010
box 0 0 192 200
use NOR3X1  NOR3X1_6
timestamp 1556798218
transform 1 0 5736 0 1 5010
box 0 0 128 200
use INVX1  INVX1_74
timestamp 1556798218
transform 1 0 5864 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_76
timestamp 1556798218
transform 1 0 5896 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_53
timestamp 1556798218
transform 1 0 5960 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_72
timestamp 1556798218
transform 1 0 6152 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_71
timestamp 1556798218
transform 1 0 6216 0 1 5010
box 0 0 64 200
use AOI22X1  AOI22X1_24
timestamp 1556798218
transform 1 0 6280 0 1 5010
box 0 0 80 200
use FILL  FILL_25_3_0
timestamp 1556798218
transform -1 0 6376 0 1 5010
box 0 0 16 200
use FILL  FILL_25_3_1
timestamp 1556798218
transform -1 0 6392 0 1 5010
box 0 0 16 200
use FILL  FILL_25_3_2
timestamp 1556798218
transform -1 0 6408 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_92
timestamp 1556798218
transform -1 0 6456 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_89
timestamp 1556798218
transform -1 0 6504 0 1 5010
box 0 0 48 200
use INVX1  INVX1_72
timestamp 1556798218
transform -1 0 6536 0 1 5010
box 0 0 32 200
use INVX1  INVX1_71
timestamp 1556798218
transform -1 0 6568 0 1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_56
timestamp 1556798218
transform -1 0 6760 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_57
timestamp 1556798218
transform -1 0 6952 0 1 5010
box 0 0 192 200
use INVX1  INVX1_75
timestamp 1556798218
transform 1 0 6952 0 1 5010
box 0 0 32 200
use NOR2X1  NOR2X1_39
timestamp 1556798218
transform -1 0 7032 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_464
timestamp 1556798218
transform 1 0 7032 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_465
timestamp 1556798218
transform -1 0 7128 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_484
timestamp 1556798218
transform -1 0 7192 0 1 5010
box 0 0 64 200
use INVX1  INVX1_543
timestamp 1556798218
transform -1 0 7224 0 1 5010
box 0 0 32 200
use AND2X2  AND2X2_69
timestamp 1556798218
transform 1 0 7224 0 1 5010
box 0 0 64 200
use AND2X2  AND2X2_15
timestamp 1556798218
transform -1 0 7352 0 1 5010
box 0 0 64 200
use INVX1  INVX1_278
timestamp 1556798218
transform 1 0 7352 0 1 5010
box 0 0 32 200
use NOR2X1  NOR2X1_102
timestamp 1556798218
transform -1 0 7432 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_175
timestamp 1556798218
transform 1 0 7432 0 1 5010
box 0 0 192 200
use INVX1  INVX1_291
timestamp 1556798218
transform 1 0 7624 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_267
timestamp 1556798218
transform 1 0 7656 0 1 5010
box 0 0 64 200
use INVX1  INVX1_290
timestamp 1556798218
transform 1 0 7720 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_265
timestamp 1556798218
transform 1 0 7752 0 1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_105
timestamp 1556798218
transform 1 0 7816 0 1 5010
box 0 0 48 200
use AOI22X1  AOI22X1_87
timestamp 1556798218
transform -1 0 7944 0 1 5010
box 0 0 80 200
use NAND2X1  NAND2X1_262
timestamp 1556798218
transform 1 0 7944 0 1 5010
box 0 0 48 200
use INVX1  INVX1_289
timestamp 1556798218
transform 1 0 7992 0 1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_43
timestamp 1556798218
transform 1 0 8024 0 1 5010
box 0 0 64 200
use BUFX2  BUFX2_136
timestamp 1556798218
transform -1 0 8136 0 1 5010
box 0 0 48 200
use FILL  FILL_26_1
timestamp 1556798218
transform 1 0 8136 0 1 5010
box 0 0 16 200
use FILL  FILL_26_2
timestamp 1556798218
transform 1 0 8152 0 1 5010
box 0 0 16 200
use INVX1  INVX1_134
timestamp 1556798218
transform 1 0 8 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_139
timestamp 1556798218
transform 1 0 40 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_130
timestamp 1556798218
transform 1 0 88 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_126
timestamp 1556798218
transform -1 0 216 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_127
timestamp 1556798218
transform -1 0 280 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_140
timestamp 1556798218
transform 1 0 280 0 -1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_47
timestamp 1556798218
transform -1 0 392 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_46
timestamp 1556798218
transform 1 0 392 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_132
timestamp 1556798218
transform 1 0 456 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_128
timestamp 1556798218
transform 1 0 488 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_138
timestamp 1556798218
transform 1 0 552 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_129
timestamp 1556798218
transform -1 0 664 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_86
timestamp 1556798218
transform 1 0 664 0 -1 5010
box 0 0 192 200
use CLKBUF1  CLKBUF1_3
timestamp 1556798218
transform 1 0 856 0 -1 5010
box 0 0 144 200
use XNOR2X1  XNOR2X1_9
timestamp 1556798218
transform 1 0 1000 0 -1 5010
box 0 0 112 200
use BUFX2  BUFX2_53
timestamp 1556798218
transform -1 0 1160 0 -1 5010
box 0 0 48 200
use INVX1  INVX1_93
timestamp 1556798218
transform -1 0 1192 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_105
timestamp 1556798218
transform 1 0 1192 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_91
timestamp 1556798218
transform 1 0 1240 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_89
timestamp 1556798218
transform 1 0 1304 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_90
timestamp 1556798218
transform -1 0 1432 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_90
timestamp 1556798218
transform -1 0 1464 0 -1 5010
box 0 0 32 200
use INVX1  INVX1_91
timestamp 1556798218
transform -1 0 1496 0 -1 5010
box 0 0 32 200
use AOI22X1  AOI22X1_30
timestamp 1556798218
transform 1 0 1496 0 -1 5010
box 0 0 80 200
use INVX1  INVX1_92
timestamp 1556798218
transform 1 0 1576 0 -1 5010
box 0 0 32 200
use CLKBUF1  CLKBUF1_7
timestamp 1556798218
transform 1 0 1608 0 -1 5010
box 0 0 144 200
use FILL  FILL_24_0_0
timestamp 1556798218
transform 1 0 1752 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_0_1
timestamp 1556798218
transform 1 0 1768 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_0_2
timestamp 1556798218
transform 1 0 1784 0 -1 5010
box 0 0 16 200
use CLKBUF1  CLKBUF1_44
timestamp 1556798218
transform 1 0 1800 0 -1 5010
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_137
timestamp 1556798218
transform 1 0 1944 0 -1 5010
box 0 0 192 200
use NAND3X1  NAND3X1_71
timestamp 1556798218
transform 1 0 2136 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_217
timestamp 1556798218
transform -1 0 2232 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_201
timestamp 1556798218
transform -1 0 2296 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_200
timestamp 1556798218
transform -1 0 2360 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_70
timestamp 1556798218
transform 1 0 2360 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_208
timestamp 1556798218
transform 1 0 2424 0 -1 5010
box 0 0 48 200
use AOI22X1  AOI22X1_66
timestamp 1556798218
transform 1 0 2472 0 -1 5010
box 0 0 80 200
use INVX1  INVX1_218
timestamp 1556798218
transform -1 0 2584 0 -1 5010
box 0 0 32 200
use BUFX2  BUFX2_55
timestamp 1556798218
transform 1 0 2584 0 -1 5010
box 0 0 48 200
use NOR2X1  NOR2X1_84
timestamp 1556798218
transform -1 0 2680 0 -1 5010
box 0 0 48 200
use AND2X2  AND2X2_59
timestamp 1556798218
transform 1 0 2680 0 -1 5010
box 0 0 64 200
use AOI22X1  AOI22X1_67
timestamp 1556798218
transform -1 0 2824 0 -1 5010
box 0 0 80 200
use OAI21X1  OAI21X1_205
timestamp 1556798218
transform -1 0 2888 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_221
timestamp 1556798218
transform -1 0 2920 0 -1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_135
timestamp 1556798218
transform 1 0 2920 0 -1 5010
box 0 0 192 200
use INVX1  INVX1_8
timestamp 1556798218
transform 1 0 3112 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_5
timestamp 1556798218
transform -1 0 3208 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_11
timestamp 1556798218
transform -1 0 3240 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_201
timestamp 1556798218
transform 1 0 3240 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_1_0
timestamp 1556798218
transform 1 0 3288 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_1_1
timestamp 1556798218
transform 1 0 3304 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_1_2
timestamp 1556798218
transform 1 0 3320 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_9
timestamp 1556798218
transform 1 0 3336 0 -1 5010
box 0 0 48 200
use INVX1  INVX1_212
timestamp 1556798218
transform 1 0 3384 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_205
timestamp 1556798218
transform 1 0 3416 0 -1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_204
timestamp 1556798218
transform -1 0 3512 0 -1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_68
timestamp 1556798218
transform -1 0 3576 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_210
timestamp 1556798218
transform 1 0 3576 0 -1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_133
timestamp 1556798218
transform -1 0 3800 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_1
timestamp 1556798218
transform -1 0 3864 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_6
timestamp 1556798218
transform -1 0 3896 0 -1 5010
box 0 0 32 200
use INVX1  INVX1_10
timestamp 1556798218
transform 1 0 3896 0 -1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1556798218
transform 1 0 3928 0 -1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_5
timestamp 1556798218
transform 1 0 4120 0 -1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_278
timestamp 1556798218
transform 1 0 4168 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_422
timestamp 1556798218
transform -1 0 4424 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_472
timestamp 1556798218
transform -1 0 4456 0 -1 5010
box 0 0 32 200
use CLKBUF1  CLKBUF1_9
timestamp 1556798218
transform -1 0 4600 0 -1 5010
box 0 0 144 200
use BUFX2  BUFX2_90
timestamp 1556798218
transform 1 0 4600 0 -1 5010
box 0 0 48 200
use AND2X2  AND2X2_118
timestamp 1556798218
transform 1 0 4648 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_10
timestamp 1556798218
transform -1 0 4760 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_2_0
timestamp 1556798218
transform -1 0 4776 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_2_1
timestamp 1556798218
transform -1 0 4792 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_2_2
timestamp 1556798218
transform -1 0 4808 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_281
timestamp 1556798218
transform -1 0 5000 0 -1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_49
timestamp 1556798218
transform -1 0 5192 0 -1 5010
box 0 0 192 200
use BUFX2  BUFX2_32
timestamp 1556798218
transform 1 0 5192 0 -1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_48
timestamp 1556798218
transform -1 0 5432 0 -1 5010
box 0 0 192 200
use NAND3X1  NAND3X1_27
timestamp 1556798218
transform 1 0 5432 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_434
timestamp 1556798218
transform -1 0 5544 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_70
timestamp 1556798218
transform -1 0 5608 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_67
timestamp 1556798218
transform -1 0 5640 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_80
timestamp 1556798218
transform 1 0 5640 0 -1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_81
timestamp 1556798218
transform 1 0 5688 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_64
timestamp 1556798218
transform 1 0 5736 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_51
timestamp 1556798218
transform -1 0 5992 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_435
timestamp 1556798218
transform -1 0 6040 0 -1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_55
timestamp 1556798218
transform 1 0 6040 0 -1 5010
box 0 0 192 200
use INVX1  INVX1_81
timestamp 1556798218
transform 1 0 6232 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_82
timestamp 1556798218
transform 1 0 6264 0 -1 5010
box 0 0 64 200
use FILL  FILL_24_3_0
timestamp 1556798218
transform 1 0 6328 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_3_1
timestamp 1556798218
transform 1 0 6344 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_3_2
timestamp 1556798218
transform 1 0 6360 0 -1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_80
timestamp 1556798218
transform 1 0 6376 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_54
timestamp 1556798218
transform 1 0 6440 0 -1 5010
box 0 0 192 200
use INVX1  INVX1_79
timestamp 1556798218
transform 1 0 6632 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_79
timestamp 1556798218
transform -1 0 6728 0 -1 5010
box 0 0 64 200
use AOI22X1  AOI22X1_26
timestamp 1556798218
transform 1 0 6728 0 -1 5010
box 0 0 80 200
use INVX1  INVX1_78
timestamp 1556798218
transform 1 0 6808 0 -1 5010
box 0 0 32 200
use NAND2X1  NAND2X1_94
timestamp 1556798218
transform 1 0 6840 0 -1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_30
timestamp 1556798218
transform -1 0 6952 0 -1 5010
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1556798218
transform 1 0 6952 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1556798218
transform 1 0 7016 0 -1 5010
box 0 0 64 200
use XNOR2X1  XNOR2X1_7
timestamp 1556798218
transform -1 0 7192 0 -1 5010
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_319
timestamp 1556798218
transform 1 0 7192 0 -1 5010
box 0 0 192 200
use INVX1  INVX1_283
timestamp 1556798218
transform 1 0 7384 0 -1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_173
timestamp 1556798218
transform -1 0 7608 0 -1 5010
box 0 0 192 200
use NAND3X1  NAND3X1_89
timestamp 1556798218
transform 1 0 7608 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_257
timestamp 1556798218
transform 1 0 7672 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_280
timestamp 1556798218
transform 1 0 7736 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_256
timestamp 1556798218
transform -1 0 7832 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_260
timestamp 1556798218
transform -1 0 7896 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_258
timestamp 1556798218
transform -1 0 7944 0 -1 5010
box 0 0 48 200
use AND2X2  AND2X2_70
timestamp 1556798218
transform -1 0 8008 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_265
timestamp 1556798218
transform 1 0 8008 0 -1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_266
timestamp 1556798218
transform -1 0 8104 0 -1 5010
box 0 0 48 200
use INVX1  INVX1_267
timestamp 1556798218
transform 1 0 8104 0 -1 5010
box 0 0 32 200
use FILL  FILL_25_1
timestamp 1556798218
transform -1 0 8152 0 -1 5010
box 0 0 16 200
use FILL  FILL_25_2
timestamp 1556798218
transform -1 0 8168 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_87
timestamp 1556798218
transform -1 0 200 0 1 4610
box 0 0 192 200
use INVX1  INVX1_137
timestamp 1556798218
transform 1 0 200 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_131
timestamp 1556798218
transform 1 0 232 0 1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_42
timestamp 1556798218
transform -1 0 376 0 1 4610
box 0 0 80 200
use INVX1  INVX1_133
timestamp 1556798218
transform -1 0 408 0 1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_89
timestamp 1556798218
transform 1 0 408 0 1 4610
box 0 0 192 200
use NAND2X1  NAND2X1_141
timestamp 1556798218
transform -1 0 648 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_142
timestamp 1556798218
transform 1 0 648 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_58
timestamp 1556798218
transform -1 0 744 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_43
timestamp 1556798218
transform -1 0 824 0 1 4610
box 0 0 80 200
use AND2X2  AND2X2_45
timestamp 1556798218
transform -1 0 888 0 1 4610
box 0 0 64 200
use INVX1  INVX1_136
timestamp 1556798218
transform -1 0 920 0 1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_368
timestamp 1556798218
transform 1 0 920 0 1 4610
box 0 0 192 200
use INVX1  INVX1_621
timestamp 1556798218
transform 1 0 1112 0 1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_243
timestamp 1556798218
transform -1 0 1192 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_62
timestamp 1556798218
transform -1 0 1384 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_92
timestamp 1556798218
transform -1 0 1448 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_104
timestamp 1556798218
transform -1 0 1496 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_108
timestamp 1556798218
transform 1 0 1496 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_107
timestamp 1556798218
transform -1 0 1592 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_45
timestamp 1556798218
transform -1 0 1640 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_31
timestamp 1556798218
transform -1 0 1720 0 1 4610
box 0 0 80 200
use FILL  FILL_23_0_0
timestamp 1556798218
transform -1 0 1736 0 1 4610
box 0 0 16 200
use FILL  FILL_23_0_1
timestamp 1556798218
transform -1 0 1752 0 1 4610
box 0 0 16 200
use FILL  FILL_23_0_2
timestamp 1556798218
transform -1 0 1768 0 1 4610
box 0 0 16 200
use AND2X2  AND2X2_38
timestamp 1556798218
transform -1 0 1832 0 1 4610
box 0 0 64 200
use INVX1  INVX1_94
timestamp 1556798218
transform -1 0 1864 0 1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_15
timestamp 1556798218
transform 1 0 1864 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_235
timestamp 1556798218
transform -1 0 2104 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_358
timestamp 1556798218
transform 1 0 2104 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_351
timestamp 1556798218
transform -1 0 2216 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_117
timestamp 1556798218
transform 1 0 2216 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_148
timestamp 1556798218
transform 1 0 2296 0 1 4610
box 0 0 48 200
use INVX1  INVX1_393
timestamp 1556798218
transform -1 0 2376 0 1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_116
timestamp 1556798218
transform 1 0 2376 0 1 4610
box 0 0 80 200
use INVX1  INVX1_394
timestamp 1556798218
transform 1 0 2456 0 1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_349
timestamp 1556798218
transform -1 0 2536 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_355
timestamp 1556798218
transform 1 0 2536 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_234
timestamp 1556798218
transform -1 0 2792 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_356
timestamp 1556798218
transform -1 0 2856 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_236
timestamp 1556798218
transform -1 0 3048 0 1 4610
box 0 0 192 200
use INVX1  INVX1_395
timestamp 1556798218
transform -1 0 3080 0 1 4610
box 0 0 32 200
use BUFX2  BUFX2_88
timestamp 1556798218
transform -1 0 3128 0 1 4610
box 0 0 48 200
use AND2X2  AND2X2_92
timestamp 1556798218
transform -1 0 3192 0 1 4610
box 0 0 64 200
use BUFX2  BUFX2_92
timestamp 1556798218
transform 1 0 3192 0 1 4610
box 0 0 48 200
use FILL  FILL_23_1_0
timestamp 1556798218
transform -1 0 3256 0 1 4610
box 0 0 16 200
use FILL  FILL_23_1_1
timestamp 1556798218
transform -1 0 3272 0 1 4610
box 0 0 16 200
use FILL  FILL_23_1_2
timestamp 1556798218
transform -1 0 3288 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_132
timestamp 1556798218
transform -1 0 3480 0 1 4610
box 0 0 192 200
use AOI21X1  AOI21X1_31
timestamp 1556798218
transform 1 0 3480 0 1 4610
box 0 0 64 200
use INVX1  INVX1_209
timestamp 1556798218
transform 1 0 3544 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_198
timestamp 1556798218
transform -1 0 3640 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_202
timestamp 1556798218
transform -1 0 3688 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_69
timestamp 1556798218
transform 1 0 3688 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_195
timestamp 1556798218
transform 1 0 3752 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_194
timestamp 1556798218
transform -1 0 3880 0 1 4610
box 0 0 64 200
use INVX1  INVX1_211
timestamp 1556798218
transform -1 0 3912 0 1 4610
box 0 0 32 200
use INVX1  INVX1_611
timestamp 1556798218
transform 1 0 3912 0 1 4610
box 0 0 32 200
use AOI21X1  AOI21X1_88
timestamp 1556798218
transform -1 0 4008 0 1 4610
box 0 0 64 200
use XNOR2X1  XNOR2X1_83
timestamp 1556798218
transform -1 0 4120 0 1 4610
box 0 0 112 200
use NAND2X1  NAND2X1_519
timestamp 1556798218
transform 1 0 4120 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_360
timestamp 1556798218
transform 1 0 4168 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_91
timestamp 1556798218
transform -1 0 4408 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_408
timestamp 1556798218
transform 1 0 4408 0 1 4610
box 0 0 48 200
use AND2X2  AND2X2_109
timestamp 1556798218
transform 1 0 4456 0 1 4610
box 0 0 64 200
use INVX1  INVX1_468
timestamp 1556798218
transform 1 0 4520 0 1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_139
timestamp 1556798218
transform 1 0 4552 0 1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_421
timestamp 1556798218
transform -1 0 4696 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_182
timestamp 1556798218
transform 1 0 4696 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_138
timestamp 1556798218
transform 1 0 4744 0 1 4610
box 0 0 80 200
use FILL  FILL_23_2_0
timestamp 1556798218
transform -1 0 4840 0 1 4610
box 0 0 16 200
use FILL  FILL_23_2_1
timestamp 1556798218
transform -1 0 4856 0 1 4610
box 0 0 16 200
use FILL  FILL_23_2_2
timestamp 1556798218
transform -1 0 4872 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_410
timestamp 1556798218
transform -1 0 4920 0 1 4610
box 0 0 48 200
use INVX1  INVX1_470
timestamp 1556798218
transform 1 0 4920 0 1 4610
box 0 0 32 200
use NAND3X1  NAND3X1_142
timestamp 1556798218
transform -1 0 5016 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_419
timestamp 1556798218
transform 1 0 5016 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_420
timestamp 1556798218
transform -1 0 5144 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_143
timestamp 1556798218
transform -1 0 5208 0 1 4610
box 0 0 64 200
use XNOR2X1  XNOR2X1_5
timestamp 1556798218
transform -1 0 5320 0 1 4610
box 0 0 112 200
use AOI21X1  AOI21X1_10
timestamp 1556798218
transform 1 0 5320 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_69
timestamp 1556798218
transform -1 0 5448 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_83
timestamp 1556798218
transform 1 0 5448 0 1 4610
box 0 0 48 200
use INVX1  INVX1_63
timestamp 1556798218
transform 1 0 5496 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_66
timestamp 1556798218
transform 1 0 5528 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_65
timestamp 1556798218
transform -1 0 5656 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_26
timestamp 1556798218
transform 1 0 5656 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_84
timestamp 1556798218
transform 1 0 5720 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_22
timestamp 1556798218
transform 1 0 5768 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_36
timestamp 1556798218
transform -1 0 5896 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_85
timestamp 1556798218
transform 1 0 5896 0 1 4610
box 0 0 48 200
use INVX1  INVX1_64
timestamp 1556798218
transform -1 0 5976 0 1 4610
box 0 0 32 200
use BUFX2  BUFX2_44
timestamp 1556798218
transform -1 0 6024 0 1 4610
box 0 0 48 200
use AND2X2  AND2X2_19
timestamp 1556798218
transform 1 0 6024 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1556798218
transform -1 0 6136 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_28
timestamp 1556798218
transform 1 0 6136 0 1 4610
box 0 0 48 200
use INVX1  INVX1_59
timestamp 1556798218
transform -1 0 6216 0 1 4610
box 0 0 32 200
use AND2X2  AND2X2_32
timestamp 1556798218
transform 1 0 6216 0 1 4610
box 0 0 64 200
use BUFX2  BUFX2_43
timestamp 1556798218
transform -1 0 6328 0 1 4610
box 0 0 48 200
use INVX1  INVX1_80
timestamp 1556798218
transform -1 0 6360 0 1 4610
box 0 0 32 200
use FILL  FILL_23_3_0
timestamp 1556798218
transform -1 0 6376 0 1 4610
box 0 0 16 200
use FILL  FILL_23_3_1
timestamp 1556798218
transform -1 0 6392 0 1 4610
box 0 0 16 200
use FILL  FILL_23_3_2
timestamp 1556798218
transform -1 0 6408 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_64
timestamp 1556798218
transform -1 0 6456 0 1 4610
box 0 0 48 200
use AND2X2  AND2X2_35
timestamp 1556798218
transform 1 0 6456 0 1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_27
timestamp 1556798218
transform 1 0 6520 0 1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_96
timestamp 1556798218
transform 1 0 6600 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_95
timestamp 1556798218
transform -1 0 6696 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_42
timestamp 1556798218
transform 1 0 6696 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_45
timestamp 1556798218
transform 1 0 6744 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_40
timestamp 1556798218
transform -1 0 6840 0 1 4610
box 0 0 48 200
use INVX1  INVX1_77
timestamp 1556798218
transform 1 0 6840 0 1 4610
box 0 0 32 200
use INVX1  INVX1_76
timestamp 1556798218
transform 1 0 6872 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_77
timestamp 1556798218
transform 1 0 6904 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_81
timestamp 1556798218
transform 1 0 6968 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_78
timestamp 1556798218
transform -1 0 7096 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_93
timestamp 1556798218
transform -1 0 7144 0 1 4610
box 0 0 48 200
use INVX1  INVX1_572
timestamp 1556798218
transform 1 0 7144 0 1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_223
timestamp 1556798218
transform -1 0 7224 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_170
timestamp 1556798218
transform 1 0 7224 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_259
timestamp 1556798218
transform 1 0 7416 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_258
timestamp 1556798218
transform -1 0 7544 0 1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_85
timestamp 1556798218
transform -1 0 7624 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_103
timestamp 1556798218
transform 1 0 7624 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_88
timestamp 1556798218
transform 1 0 7672 0 1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_84
timestamp 1556798218
transform 1 0 7736 0 1 4610
box 0 0 80 200
use INVX1  INVX1_281
timestamp 1556798218
transform -1 0 7848 0 1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_259
timestamp 1556798218
transform -1 0 7896 0 1 4610
box 0 0 48 200
use INVX1  INVX1_279
timestamp 1556798218
transform -1 0 7928 0 1 4610
box 0 0 32 200
use INVX1  INVX1_282
timestamp 1556798218
transform -1 0 7960 0 1 4610
box 0 0 32 200
use AOI21X1  AOI21X1_41
timestamp 1556798218
transform -1 0 8024 0 1 4610
box 0 0 64 200
use XNOR2X1  XNOR2X1_36
timestamp 1556798218
transform -1 0 8136 0 1 4610
box 0 0 112 200
use FILL  FILL_24_1
timestamp 1556798218
transform 1 0 8136 0 1 4610
box 0 0 16 200
use FILL  FILL_24_2
timestamp 1556798218
transform 1 0 8152 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_346
timestamp 1556798218
transform -1 0 200 0 -1 4610
box 0 0 192 200
use AND2X2  AND2X2_43
timestamp 1556798218
transform 1 0 200 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_176
timestamp 1556798218
transform -1 0 328 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_587
timestamp 1556798218
transform -1 0 360 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_521
timestamp 1556798218
transform 1 0 360 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_522
timestamp 1556798218
transform 1 0 424 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_177
timestamp 1556798218
transform -1 0 552 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_233
timestamp 1556798218
transform 1 0 552 0 -1 4610
box 0 0 48 200
use INVX1  INVX1_586
timestamp 1556798218
transform -1 0 632 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_349
timestamp 1556798218
transform 1 0 632 0 -1 4610
box 0 0 192 200
use AOI21X1  AOI21X1_90
timestamp 1556798218
transform 1 0 824 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_555
timestamp 1556798218
transform -1 0 952 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_623
timestamp 1556798218
transform 1 0 952 0 -1 4610
box 0 0 32 200
use INVX1  INVX1_625
timestamp 1556798218
transform -1 0 1016 0 -1 4610
box 0 0 32 200
use NAND3X1  NAND3X1_187
timestamp 1556798218
transform 1 0 1016 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_369
timestamp 1556798218
transform 1 0 1080 0 -1 4610
box 0 0 192 200
use AND2X2  AND2X2_36
timestamp 1556798218
transform 1 0 1272 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_366
timestamp 1556798218
transform -1 0 1528 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_94
timestamp 1556798218
transform 1 0 1528 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_95
timestamp 1556798218
transform -1 0 1624 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_63
timestamp 1556798218
transform 1 0 1624 0 -1 4610
box 0 0 192 200
use FILL  FILL_22_0_0
timestamp 1556798218
transform -1 0 1832 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_1
timestamp 1556798218
transform -1 0 1848 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_2
timestamp 1556798218
transform -1 0 1864 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_201
timestamp 1556798218
transform -1 0 2056 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_396
timestamp 1556798218
transform 1 0 2056 0 -1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_350
timestamp 1556798218
transform 1 0 2088 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_237
timestamp 1556798218
transform -1 0 2328 0 -1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_121
timestamp 1556798218
transform -1 0 2392 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_354
timestamp 1556798218
transform 1 0 2392 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_120
timestamp 1556798218
transform -1 0 2520 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_353
timestamp 1556798218
transform 1 0 2520 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_392
timestamp 1556798218
transform 1 0 2584 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_357
timestamp 1556798218
transform 1 0 2616 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_348
timestamp 1556798218
transform -1 0 2728 0 -1 4610
box 0 0 48 200
use INVX1  INVX1_391
timestamp 1556798218
transform -1 0 2760 0 -1 4610
box 0 0 32 200
use AOI21X1  AOI21X1_57
timestamp 1556798218
transform -1 0 2824 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_347
timestamp 1556798218
transform -1 0 2872 0 -1 4610
box 0 0 48 200
use XNOR2X1  XNOR2X1_52
timestamp 1556798218
transform 1 0 2872 0 -1 4610
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_197
timestamp 1556798218
transform 1 0 2984 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_2
timestamp 1556798218
transform 1 0 3176 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1556798218
transform 1 0 3240 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_1_0
timestamp 1556798218
transform 1 0 3304 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_1
timestamp 1556798218
transform 1 0 3320 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_2
timestamp 1556798218
transform 1 0 3336 0 -1 4610
box 0 0 16 200
use INVX1  INVX1_607
timestamp 1556798218
transform 1 0 3352 0 -1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_239
timestamp 1556798218
transform -1 0 3432 0 -1 4610
box 0 0 48 200
use XNOR2X1  XNOR2X1_26
timestamp 1556798218
transform 1 0 3432 0 -1 4610
box 0 0 112 200
use INVX1  INVX1_208
timestamp 1556798218
transform -1 0 3576 0 -1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_81
timestamp 1556798218
transform 1 0 3576 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_183
timestamp 1556798218
transform -1 0 3688 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_543
timestamp 1556798218
transform -1 0 3752 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_539
timestamp 1556798218
transform -1 0 3816 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_13
timestamp 1556798218
transform 1 0 3816 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_540
timestamp 1556798218
transform -1 0 3912 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_518
timestamp 1556798218
transform -1 0 3960 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_182
timestamp 1556798218
transform 1 0 3960 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_541
timestamp 1556798218
transform 1 0 4024 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_608
timestamp 1556798218
transform -1 0 4120 0 -1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_178
timestamp 1556798218
transform 1 0 4120 0 -1 4610
box 0 0 80 200
use INVX1  INVX1_610
timestamp 1556798218
transform -1 0 4232 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_544
timestamp 1556798218
transform -1 0 4296 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_613
timestamp 1556798218
transform -1 0 4328 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_359
timestamp 1556798218
transform 1 0 4328 0 -1 4610
box 0 0 192 200
use XNOR2X1  XNOR2X1_63
timestamp 1556798218
transform -1 0 4632 0 -1 4610
box 0 0 112 200
use NAND2X1  NAND2X1_412
timestamp 1556798218
transform 1 0 4632 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_411
timestamp 1556798218
transform -1 0 4728 0 -1 4610
box 0 0 48 200
use INVX1  INVX1_471
timestamp 1556798218
transform 1 0 4728 0 -1 4610
box 0 0 32 200
use INVX1  INVX1_12
timestamp 1556798218
transform 1 0 4760 0 -1 4610
box 0 0 32 200
use FILL  FILL_22_2_0
timestamp 1556798218
transform -1 0 4808 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_1
timestamp 1556798218
transform -1 0 4824 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_2
timestamp 1556798218
transform -1 0 4840 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_280
timestamp 1556798218
transform -1 0 5032 0 -1 4610
box 0 0 192 200
use AOI21X1  AOI21X1_68
timestamp 1556798218
transform 1 0 5032 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_469
timestamp 1556798218
transform 1 0 5096 0 -1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_409
timestamp 1556798218
transform 1 0 5128 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_423
timestamp 1556798218
transform 1 0 5176 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_181
timestamp 1556798218
transform 1 0 5240 0 -1 4610
box 0 0 48 200
use INVX1  INVX1_467
timestamp 1556798218
transform -1 0 5320 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_46
timestamp 1556798218
transform 1 0 5320 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_68
timestamp 1556798218
transform 1 0 5512 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_82
timestamp 1556798218
transform -1 0 5624 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_67
timestamp 1556798218
transform -1 0 5688 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_62
timestamp 1556798218
transform 1 0 5688 0 -1 4610
box 0 0 32 200
use INVX1  INVX1_65
timestamp 1556798218
transform 1 0 5720 0 -1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_23
timestamp 1556798218
transform -1 0 5832 0 -1 4610
box 0 0 80 200
use BUFX2  BUFX2_62
timestamp 1556798218
transform 1 0 5832 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_86
timestamp 1556798218
transform 1 0 5880 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_317
timestamp 1556798218
transform -1 0 6120 0 -1 4610
box 0 0 192 200
use NAND2X1  NAND2X1_75
timestamp 1556798218
transform -1 0 6168 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_61
timestamp 1556798218
transform 1 0 6168 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_42
timestamp 1556798218
transform 1 0 6232 0 -1 4610
box 0 0 192 200
use FILL  FILL_22_3_0
timestamp 1556798218
transform 1 0 6424 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_3_1
timestamp 1556798218
transform 1 0 6440 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_3_2
timestamp 1556798218
transform 1 0 6456 0 -1 4610
box 0 0 16 200
use AOI22X1  AOI22X1_21
timestamp 1556798218
transform 1 0 6472 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_60
timestamp 1556798218
transform -1 0 6616 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_34
timestamp 1556798218
transform 1 0 6616 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_63
timestamp 1556798218
transform -1 0 6728 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_60
timestamp 1556798218
transform -1 0 6760 0 -1 4610
box 0 0 32 200
use INVX1  INVX1_55
timestamp 1556798218
transform -1 0 6792 0 -1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_20
timestamp 1556798218
transform 1 0 6792 0 -1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_77
timestamp 1556798218
transform -1 0 6920 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_43
timestamp 1556798218
transform 1 0 6920 0 -1 4610
box 0 0 192 200
use AOI21X1  AOI21X1_83
timestamp 1556798218
transform 1 0 7112 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_340
timestamp 1556798218
transform 1 0 7176 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_513
timestamp 1556798218
transform -1 0 7432 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_490
timestamp 1556798218
transform -1 0 7480 0 -1 4610
box 0 0 48 200
use AND2X2  AND2X2_17
timestamp 1556798218
transform 1 0 7480 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_257
timestamp 1556798218
transform 1 0 7544 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_261
timestamp 1556798218
transform 1 0 7592 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_260
timestamp 1556798218
transform -1 0 7688 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_261
timestamp 1556798218
transform -1 0 7752 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_171
timestamp 1556798218
transform -1 0 7944 0 -1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_172
timestamp 1556798218
transform -1 0 8136 0 -1 4610
box 0 0 192 200
use FILL  FILL_23_1
timestamp 1556798218
transform -1 0 8152 0 -1 4610
box 0 0 16 200
use FILL  FILL_23_2
timestamp 1556798218
transform -1 0 8168 0 -1 4610
box 0 0 16 200
use INVX1  INVX1_591
timestamp 1556798218
transform -1 0 40 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_524
timestamp 1556798218
transform 1 0 40 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_523
timestamp 1556798218
transform -1 0 168 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_234
timestamp 1556798218
transform -1 0 216 0 1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_172
timestamp 1556798218
transform 1 0 216 0 1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_504
timestamp 1556798218
transform -1 0 344 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_505
timestamp 1556798218
transform 1 0 344 0 1 4210
box 0 0 48 200
use INVX1  INVX1_589
timestamp 1556798218
transform -1 0 424 0 1 4210
box 0 0 32 200
use INVX1  INVX1_590
timestamp 1556798218
transform -1 0 456 0 1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_85
timestamp 1556798218
transform 1 0 456 0 1 4210
box 0 0 64 200
use XNOR2X1  XNOR2X1_80
timestamp 1556798218
transform -1 0 632 0 1 4210
box 0 0 112 200
use OAI21X1  OAI21X1_525
timestamp 1556798218
transform -1 0 696 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_503
timestamp 1556798218
transform -1 0 744 0 1 4210
box 0 0 48 200
use INVX1  INVX1_588
timestamp 1556798218
transform -1 0 776 0 1 4210
box 0 0 32 200
use BUFX2  BUFX2_12
timestamp 1556798218
transform -1 0 824 0 1 4210
box 0 0 48 200
use XNOR2X1  XNOR2X1_85
timestamp 1556798218
transform -1 0 936 0 1 4210
box 0 0 112 200
use NAND2X1  NAND2X1_528
timestamp 1556798218
transform 1 0 936 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_551
timestamp 1556798218
transform -1 0 1048 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_552
timestamp 1556798218
transform -1 0 1112 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_186
timestamp 1556798218
transform 1 0 1112 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_182
timestamp 1556798218
transform -1 0 1256 0 1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_529
timestamp 1556798218
transform -1 0 1304 0 1 4210
box 0 0 48 200
use INVX1  INVX1_622
timestamp 1556798218
transform -1 0 1336 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_553
timestamp 1556798218
transform 1 0 1336 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_527
timestamp 1556798218
transform 1 0 1400 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_554
timestamp 1556798218
transform 1 0 1448 0 1 4210
box 0 0 64 200
use INVX1  INVX1_332
timestamp 1556798218
transform 1 0 1512 0 1 4210
box 0 0 32 200
use AND2X2  AND2X2_21
timestamp 1556798218
transform 1 0 1544 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_302
timestamp 1556798218
transform 1 0 1608 0 1 4210
box 0 0 64 200
use FILL  FILL_21_0_0
timestamp 1556798218
transform 1 0 1672 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_1
timestamp 1556798218
transform 1 0 1688 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_2
timestamp 1556798218
transform 1 0 1704 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_198
timestamp 1556798218
transform 1 0 1720 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_301
timestamp 1556798218
transform -1 0 1976 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_102
timestamp 1556798218
transform -1 0 2040 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_103
timestamp 1556798218
transform -1 0 2104 0 1 4210
box 0 0 64 200
use INVX1  INVX1_327
timestamp 1556798218
transform 1 0 2104 0 1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_117
timestamp 1556798218
transform -1 0 2184 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_300
timestamp 1556798218
transform 1 0 2184 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_299
timestamp 1556798218
transform 1 0 2248 0 1 4210
box 0 0 64 200
use INVX1  INVX1_329
timestamp 1556798218
transform 1 0 2312 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_303
timestamp 1556798218
transform 1 0 2344 0 1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_48
timestamp 1556798218
transform 1 0 2408 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_200
timestamp 1556798218
transform -1 0 2664 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_294
timestamp 1556798218
transform -1 0 2728 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_292
timestamp 1556798218
transform -1 0 2776 0 1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_147
timestamp 1556798218
transform 1 0 2776 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_297
timestamp 1556798218
transform 1 0 2824 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_101
timestamp 1556798218
transform -1 0 2952 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_115
timestamp 1556798218
transform 1 0 2952 0 1 4210
box 0 0 48 200
use INVX1  INVX1_390
timestamp 1556798218
transform -1 0 3032 0 1 4210
box 0 0 32 200
use INVX1  INVX1_320
timestamp 1556798218
transform -1 0 3064 0 1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_192
timestamp 1556798218
transform -1 0 3256 0 1 4210
box 0 0 192 200
use BUFX2  BUFX2_30
timestamp 1556798218
transform -1 0 3304 0 1 4210
box 0 0 48 200
use FILL  FILL_21_1_0
timestamp 1556798218
transform -1 0 3320 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_1
timestamp 1556798218
transform -1 0 3336 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_2
timestamp 1556798218
transform -1 0 3352 0 1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_7
timestamp 1556798218
transform -1 0 3416 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_6
timestamp 1556798218
transform 1 0 3416 0 1 4210
box 0 0 64 200
use BUFX2  BUFX2_9
timestamp 1556798218
transform 1 0 3480 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_361
timestamp 1556798218
transform -1 0 3720 0 1 4210
box 0 0 192 200
use INVX1  INVX1_609
timestamp 1556798218
transform 1 0 3720 0 1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_240
timestamp 1556798218
transform 1 0 3752 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_520
timestamp 1556798218
transform 1 0 3800 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_521
timestamp 1556798218
transform -1 0 3896 0 1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_179
timestamp 1556798218
transform 1 0 3896 0 1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_517
timestamp 1556798218
transform 1 0 3976 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_542
timestamp 1556798218
transform 1 0 4024 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_358
timestamp 1556798218
transform -1 0 4280 0 1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_9
timestamp 1556798218
transform 1 0 4280 0 1 4210
box 0 0 64 200
use INVX1  INVX1_3
timestamp 1556798218
transform -1 0 4376 0 1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_1
timestamp 1556798218
transform -1 0 4440 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1556798218
transform 1 0 4440 0 1 4210
box 0 0 64 200
use INVX1  INVX1_473
timestamp 1556798218
transform 1 0 4504 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_424
timestamp 1556798218
transform 1 0 4536 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_279
timestamp 1556798218
transform 1 0 4600 0 1 4210
box 0 0 192 200
use FILL  FILL_21_2_0
timestamp 1556798218
transform 1 0 4792 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_1
timestamp 1556798218
transform 1 0 4808 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_2
timestamp 1556798218
transform 1 0 4824 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_6
timestamp 1556798218
transform 1 0 4840 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_10
timestamp 1556798218
transform -1 0 4968 0 1 4210
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1556798218
transform 1 0 4968 0 1 4210
box 0 0 64 200
use XOR2X1  XOR2X1_1
timestamp 1556798218
transform -1 0 5144 0 1 4210
box 0 0 112 200
use NAND2X1  NAND2X1_60
timestamp 1556798218
transform -1 0 5192 0 1 4210
box 0 0 48 200
use BUFX2  BUFX2_65
timestamp 1556798218
transform -1 0 5240 0 1 4210
box 0 0 48 200
use AND2X2  AND2X2_33
timestamp 1556798218
transform 1 0 5240 0 1 4210
box 0 0 64 200
use INVX1  INVX1_66
timestamp 1556798218
transform 1 0 5304 0 1 4210
box 0 0 32 200
use AND2X2  AND2X2_28
timestamp 1556798218
transform 1 0 5336 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_314
timestamp 1556798218
transform 1 0 5400 0 1 4210
box 0 0 192 200
use AND2X2  AND2X2_121
timestamp 1556798218
transform 1 0 5592 0 1 4210
box 0 0 64 200
use INVX1  INVX1_535
timestamp 1556798218
transform 1 0 5656 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_476
timestamp 1556798218
transform 1 0 5688 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_475
timestamp 1556798218
transform -1 0 5816 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_157
timestamp 1556798218
transform 1 0 5816 0 1 4210
box 0 0 80 200
use NOR2X1  NOR2X1_206
timestamp 1556798218
transform -1 0 5944 0 1 4210
box 0 0 48 200
use INVX1  INVX1_532
timestamp 1556798218
transform 1 0 5944 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_473
timestamp 1556798218
transform 1 0 5976 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_474
timestamp 1556798218
transform -1 0 6104 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_161
timestamp 1556798218
transform -1 0 6168 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_160
timestamp 1556798218
transform 1 0 6168 0 1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_77
timestamp 1556798218
transform 1 0 6232 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_477
timestamp 1556798218
transform 1 0 6296 0 1 4210
box 0 0 64 200
use FILL  FILL_21_3_0
timestamp 1556798218
transform -1 0 6376 0 1 4210
box 0 0 16 200
use FILL  FILL_21_3_1
timestamp 1556798218
transform -1 0 6392 0 1 4210
box 0 0 16 200
use FILL  FILL_21_3_2
timestamp 1556798218
transform -1 0 6408 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_457
timestamp 1556798218
transform -1 0 6456 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_79
timestamp 1556798218
transform -1 0 6504 0 1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_205
timestamp 1556798218
transform 1 0 6504 0 1 4210
box 0 0 48 200
use INVX1  INVX1_530
timestamp 1556798218
transform -1 0 6584 0 1 4210
box 0 0 32 200
use INVX1  INVX1_58
timestamp 1556798218
transform 1 0 6584 0 1 4210
box 0 0 32 200
use INVX1  INVX1_57
timestamp 1556798218
transform 1 0 6616 0 1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_9
timestamp 1556798218
transform -1 0 6712 0 1 4210
box 0 0 64 200
use XNOR2X1  XNOR2X1_4
timestamp 1556798218
transform 1 0 6712 0 1 4210
box 0 0 112 200
use NAND3X1  NAND3X1_24
timestamp 1556798218
transform 1 0 6824 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1556798218
transform 1 0 6888 0 1 4210
box 0 0 64 200
use INVX1  INVX1_56
timestamp 1556798218
transform 1 0 6952 0 1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_341
timestamp 1556798218
transform -1 0 7176 0 1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_172
timestamp 1556798218
transform -1 0 7240 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_173
timestamp 1556798218
transform -1 0 7304 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_510
timestamp 1556798218
transform 1 0 7304 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_509
timestamp 1556798218
transform 1 0 7368 0 1 4210
box 0 0 64 200
use INVX1  INVX1_574
timestamp 1556798218
transform -1 0 7464 0 1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_491
timestamp 1556798218
transform 1 0 7464 0 1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_168
timestamp 1556798218
transform -1 0 7592 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_514
timestamp 1556798218
transform -1 0 7656 0 1 4210
box 0 0 64 200
use INVX1  INVX1_578
timestamp 1556798218
transform -1 0 7688 0 1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_251
timestamp 1556798218
transform -1 0 7736 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_250
timestamp 1556798218
transform -1 0 7784 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_249
timestamp 1556798218
transform -1 0 7848 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_339
timestamp 1556798218
transform 1 0 7848 0 1 4210
box 0 0 192 200
use BUFX2  BUFX2_57
timestamp 1556798218
transform -1 0 8088 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_234
timestamp 1556798218
transform -1 0 8136 0 1 4210
box 0 0 48 200
use FILL  FILL_22_1
timestamp 1556798218
transform 1 0 8136 0 1 4210
box 0 0 16 200
use FILL  FILL_22_2
timestamp 1556798218
transform 1 0 8152 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_526
timestamp 1556798218
transform 1 0 8 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_502
timestamp 1556798218
transform -1 0 120 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_173
timestamp 1556798218
transform -1 0 200 0 -1 4210
box 0 0 80 200
use AND2X2  AND2X2_135
timestamp 1556798218
transform -1 0 264 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_506
timestamp 1556798218
transform -1 0 312 0 -1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_348
timestamp 1556798218
transform -1 0 504 0 -1 4210
box 0 0 192 200
use BUFX2  BUFX2_26
timestamp 1556798218
transform -1 0 552 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_125
timestamp 1556798218
transform 1 0 552 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_334
timestamp 1556798218
transform -1 0 632 0 -1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_105
timestamp 1556798218
transform 1 0 632 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_205
timestamp 1556798218
transform 1 0 696 0 -1 4210
box 0 0 192 200
use INVX1  INVX1_624
timestamp 1556798218
transform 1 0 888 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_530
timestamp 1556798218
transform 1 0 920 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_531
timestamp 1556798218
transform -1 0 1016 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_244
timestamp 1556798218
transform 1 0 1016 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_183
timestamp 1556798218
transform 1 0 1064 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_556
timestamp 1556798218
transform -1 0 1208 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_627
timestamp 1556798218
transform -1 0 1240 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_367
timestamp 1556798218
transform -1 0 1432 0 -1 4210
box 0 0 192 200
use AND2X2  AND2X2_77
timestamp 1556798218
transform 1 0 1432 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_296
timestamp 1556798218
transform 1 0 1496 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_300
timestamp 1556798218
transform 1 0 1544 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_299
timestamp 1556798218
transform 1 0 1592 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_99
timestamp 1556798218
transform 1 0 1640 0 -1 4210
box 0 0 80 200
use NOR2X1  NOR2X1_118
timestamp 1556798218
transform 1 0 1720 0 -1 4210
box 0 0 48 200
use FILL  FILL_20_0_0
timestamp 1556798218
transform 1 0 1768 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_1
timestamp 1556798218
transform 1 0 1784 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_2
timestamp 1556798218
transform 1 0 1800 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_328
timestamp 1556798218
transform 1 0 1816 0 -1 4210
box 0 0 32 200
use AOI22X1  AOI22X1_98
timestamp 1556798218
transform 1 0 1848 0 -1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_298
timestamp 1556798218
transform 1 0 1928 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_331
timestamp 1556798218
transform -1 0 2008 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_330
timestamp 1556798218
transform -1 0 2040 0 -1 4210
box 0 0 32 200
use XNOR2X1  XNOR2X1_43
timestamp 1556798218
transform 1 0 2040 0 -1 4210
box 0 0 112 200
use NAND2X1  NAND2X1_297
timestamp 1556798218
transform -1 0 2200 0 -1 4210
box 0 0 48 200
use BUFX2  BUFX2_20
timestamp 1556798218
transform -1 0 2248 0 -1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_194
timestamp 1556798218
transform 1 0 2248 0 -1 4210
box 0 0 192 200
use BUFX2  BUFX2_19
timestamp 1556798218
transform 1 0 2440 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_323
timestamp 1556798218
transform 1 0 2488 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_321
timestamp 1556798218
transform 1 0 2520 0 -1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_100
timestamp 1556798218
transform -1 0 2616 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_293
timestamp 1556798218
transform 1 0 2616 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_317
timestamp 1556798218
transform 1 0 2680 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_322
timestamp 1556798218
transform -1 0 2744 0 -1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_98
timestamp 1556798218
transform -1 0 2808 0 -1 4210
box 0 0 64 200
use XNOR2X1  XNOR2X1_41
timestamp 1556798218
transform 1 0 2808 0 -1 4210
box 0 0 112 200
use NAND3X1  NAND3X1_99
timestamp 1556798218
transform -1 0 2984 0 -1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_46
timestamp 1556798218
transform 1 0 2984 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_113
timestamp 1556798218
transform 1 0 3048 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_313
timestamp 1556798218
transform -1 0 3128 0 -1 4210
box 0 0 32 200
use BUFX2  BUFX2_21
timestamp 1556798218
transform 1 0 3128 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_8
timestamp 1556798218
transform 1 0 3176 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_16
timestamp 1556798218
transform 1 0 3224 0 -1 4210
box 0 0 48 200
use FILL  FILL_20_1_0
timestamp 1556798218
transform 1 0 3272 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_1
timestamp 1556798218
transform 1 0 3288 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_2
timestamp 1556798218
transform 1 0 3304 0 -1 4210
box 0 0 16 200
use BUFX2  BUFX2_11
timestamp 1556798218
transform 1 0 3320 0 -1 4210
box 0 0 48 200
use XNOR2X1  XNOR2X1_40
timestamp 1556798218
transform -1 0 3480 0 -1 4210
box 0 0 112 200
use INVX1  INVX1_309
timestamp 1556798218
transform -1 0 3512 0 -1 4210
box 0 0 32 200
use CLKBUF1  CLKBUF1_40
timestamp 1556798218
transform -1 0 3656 0 -1 4210
box 0 0 144 200
use BUFX2  BUFX2_2
timestamp 1556798218
transform -1 0 3704 0 -1 4210
box 0 0 48 200
use AND2X2  AND2X2_138
timestamp 1556798218
transform 1 0 3704 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_612
timestamp 1556798218
transform 1 0 3768 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_7
timestamp 1556798218
transform 1 0 3800 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_11
timestamp 1556798218
transform -1 0 3928 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_4
timestamp 1556798218
transform 1 0 3928 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_23
timestamp 1556798218
transform 1 0 3992 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_24
timestamp 1556798218
transform -1 0 4088 0 -1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1556798218
transform 1 0 4088 0 -1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_26
timestamp 1556798218
transform 1 0 4280 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_12
timestamp 1556798218
transform 1 0 4328 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_2
timestamp 1556798218
transform -1 0 4424 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_4
timestamp 1556798218
transform 1 0 4424 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_10
timestamp 1556798218
transform -1 0 4504 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_27
timestamp 1556798218
transform -1 0 4552 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_8
timestamp 1556798218
transform 1 0 4552 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1556798218
transform -1 0 4744 0 -1 4210
box 0 0 128 200
use NOR2X1  NOR2X1_15
timestamp 1556798218
transform -1 0 4792 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_5
timestamp 1556798218
transform -1 0 4824 0 -1 4210
box 0 0 32 200
use FILL  FILL_20_2_0
timestamp 1556798218
transform 1 0 4824 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_1
timestamp 1556798218
transform 1 0 4840 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_2
timestamp 1556798218
transform 1 0 4856 0 -1 4210
box 0 0 16 200
use XNOR2X1  XNOR2X1_1
timestamp 1556798218
transform 1 0 4872 0 -1 4210
box 0 0 112 200
use AOI21X1  AOI21X1_6
timestamp 1556798218
transform 1 0 4984 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1556798218
transform -1 0 5112 0 -1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_5
timestamp 1556798218
transform -1 0 5176 0 -1 4210
box 0 0 64 200
use OR2X2  OR2X2_3
timestamp 1556798218
transform -1 0 5240 0 -1 4210
box 0 0 64 200
use AND2X2  AND2X2_26
timestamp 1556798218
transform -1 0 5304 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_38
timestamp 1556798218
transform 1 0 5304 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_26
timestamp 1556798218
transform 1 0 5336 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_27
timestamp 1556798218
transform 1 0 5384 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_15
timestamp 1556798218
transform 1 0 5432 0 -1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_456
timestamp 1556798218
transform 1 0 5512 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_460
timestamp 1556798218
transform 1 0 5560 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_459
timestamp 1556798218
transform -1 0 5656 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_534
timestamp 1556798218
transform 1 0 5656 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_458
timestamp 1556798218
transform 1 0 5688 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_531
timestamp 1556798218
transform 1 0 5736 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_533
timestamp 1556798218
transform 1 0 5768 0 -1 4210
box 0 0 32 200
use AOI22X1  AOI22X1_156
timestamp 1556798218
transform -1 0 5880 0 -1 4210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_316
timestamp 1556798218
transform -1 0 6072 0 -1 4210
box 0 0 192 200
use XNOR2X1  XNOR2X1_72
timestamp 1556798218
transform 1 0 6072 0 -1 4210
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_44
timestamp 1556798218
transform -1 0 6376 0 -1 4210
box 0 0 192 200
use FILL  FILL_20_3_0
timestamp 1556798218
transform -1 0 6392 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_1
timestamp 1556798218
transform -1 0 6408 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_2
timestamp 1556798218
transform -1 0 6424 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_78
timestamp 1556798218
transform -1 0 6472 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_76
timestamp 1556798218
transform 1 0 6472 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_62
timestamp 1556798218
transform 1 0 6520 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_33
timestamp 1556798218
transform 1 0 6584 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_54
timestamp 1556798218
transform -1 0 6664 0 -1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_25
timestamp 1556798218
transform 1 0 6664 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_59
timestamp 1556798218
transform 1 0 6728 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_45
timestamp 1556798218
transform 1 0 6792 0 -1 4210
box 0 0 192 200
use XNOR2X1  XNOR2X1_78
timestamp 1556798218
transform 1 0 6984 0 -1 4210
box 0 0 112 200
use INVX1  INVX1_575
timestamp 1556798218
transform 1 0 7096 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_224
timestamp 1556798218
transform -1 0 7176 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_169
timestamp 1556798218
transform 1 0 7176 0 -1 4210
box 0 0 80 200
use INVX1  INVX1_573
timestamp 1556798218
transform 1 0 7256 0 -1 4210
box 0 0 32 200
use INVX1  INVX1_576
timestamp 1556798218
transform -1 0 7320 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_511
timestamp 1556798218
transform -1 0 7384 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_493
timestamp 1556798218
transform 1 0 7384 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_492
timestamp 1556798218
transform -1 0 7480 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_264
timestamp 1556798218
transform 1 0 7480 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_98
timestamp 1556798218
transform -1 0 7560 0 -1 4210
box 0 0 48 200
use BUFX2  BUFX2_58
timestamp 1556798218
transform -1 0 7608 0 -1 4210
box 0 0 48 200
use BUFX2  BUFX2_59
timestamp 1556798218
transform 1 0 7608 0 -1 4210
box 0 0 48 200
use BUFX2  BUFX2_60
timestamp 1556798218
transform 1 0 7656 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_265
timestamp 1556798218
transform 1 0 7704 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_246
timestamp 1556798218
transform -1 0 7784 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_244
timestamp 1556798218
transform 1 0 7784 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_85
timestamp 1556798218
transform -1 0 7912 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_247
timestamp 1556798218
transform -1 0 7976 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_247
timestamp 1556798218
transform -1 0 8024 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_266
timestamp 1556798218
transform -1 0 8056 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_233
timestamp 1556798218
transform 1 0 8056 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_93
timestamp 1556798218
transform 1 0 8104 0 -1 4210
box 0 0 48 200
use FILL  FILL_21_1
timestamp 1556798218
transform -1 0 8168 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_592
timestamp 1556798218
transform -1 0 40 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_347
timestamp 1556798218
transform 1 0 40 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_304
timestamp 1556798218
transform 1 0 232 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_204
timestamp 1556798218
transform -1 0 472 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_499
timestamp 1556798218
transform -1 0 520 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_49
timestamp 1556798218
transform 1 0 520 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_309
timestamp 1556798218
transform -1 0 648 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_104
timestamp 1556798218
transform 1 0 648 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_306
timestamp 1556798218
transform 1 0 712 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_305
timestamp 1556798218
transform -1 0 840 0 1 3810
box 0 0 64 200
use INVX1  INVX1_336
timestamp 1556798218
transform -1 0 872 0 1 3810
box 0 0 32 200
use INVX1  INVX1_337
timestamp 1556798218
transform -1 0 904 0 1 3810
box 0 0 32 200
use XNOR2X1  XNOR2X1_44
timestamp 1556798218
transform -1 0 1016 0 1 3810
box 0 0 112 200
use NAND2X1  NAND2X1_307
timestamp 1556798218
transform 1 0 1016 0 1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_308
timestamp 1556798218
transform -1 0 1112 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_22
timestamp 1556798218
transform -1 0 1160 0 1 3810
box 0 0 48 200
use AND2X2  AND2X2_140
timestamp 1556798218
transform -1 0 1224 0 1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_8
timestamp 1556798218
transform 1 0 1224 0 1 3810
box 0 0 128 200
use INVX1  INVX1_626
timestamp 1556798218
transform 1 0 1352 0 1 3810
box 0 0 32 200
use BUFX2  BUFX2_10
timestamp 1556798218
transform -1 0 1432 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_58
timestamp 1556798218
transform 1 0 1432 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_86
timestamp 1556798218
transform -1 0 1688 0 1 3810
box 0 0 64 200
use INVX1  INVX1_87
timestamp 1556798218
transform -1 0 1720 0 1 3810
box 0 0 32 200
use FILL  FILL_19_0_0
timestamp 1556798218
transform -1 0 1736 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1556798218
transform -1 0 1752 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_2
timestamp 1556798218
transform -1 0 1768 0 1 3810
box 0 0 16 200
use AND2X2  AND2X2_37
timestamp 1556798218
transform -1 0 1832 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_99
timestamp 1556798218
transform 1 0 1832 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_228
timestamp 1556798218
transform -1 0 1928 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_304
timestamp 1556798218
transform -1 0 1992 0 1 3810
box 0 0 64 200
use INVX1  INVX1_333
timestamp 1556798218
transform -1 0 2024 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_195
timestamp 1556798218
transform 1 0 2024 0 1 3810
box 0 0 192 200
use INVX1  INVX1_326
timestamp 1556798218
transform 1 0 2216 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_298
timestamp 1556798218
transform 1 0 2248 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_268
timestamp 1556798218
transform -1 0 2360 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_296
timestamp 1556798218
transform 1 0 2360 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_97
timestamp 1556798218
transform -1 0 2504 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_295
timestamp 1556798218
transform -1 0 2568 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_116
timestamp 1556798218
transform -1 0 2616 0 1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_96
timestamp 1556798218
transform -1 0 2696 0 1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_293
timestamp 1556798218
transform -1 0 2744 0 1 3810
box 0 0 48 200
use INVX1  INVX1_324
timestamp 1556798218
transform 1 0 2744 0 1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_47
timestamp 1556798218
transform 1 0 2776 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_196
timestamp 1556798218
transform -1 0 3032 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_291
timestamp 1556798218
transform 1 0 3032 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_193
timestamp 1556798218
transform 1 0 3096 0 1 3810
box 0 0 192 200
use FILL  FILL_19_1_0
timestamp 1556798218
transform 1 0 3288 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1556798218
transform 1 0 3304 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_2
timestamp 1556798218
transform 1 0 3320 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_281
timestamp 1556798218
transform 1 0 3336 0 1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_92
timestamp 1556798218
transform -1 0 3464 0 1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_112
timestamp 1556798218
transform -1 0 3512 0 1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_282
timestamp 1556798218
transform 1 0 3512 0 1 3810
box 0 0 48 200
use AND2X2  AND2X2_74
timestamp 1556798218
transform 1 0 3560 0 1 3810
box 0 0 64 200
use INVX1  INVX1_311
timestamp 1556798218
transform 1 0 3624 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_283
timestamp 1556798218
transform 1 0 3656 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_282
timestamp 1556798218
transform 1 0 3720 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_93
timestamp 1556798218
transform 1 0 3784 0 1 3810
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_186
timestamp 1556798218
transform -1 0 4056 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_285
timestamp 1556798218
transform -1 0 4120 0 1 3810
box 0 0 64 200
use INVX1  INVX1_312
timestamp 1556798218
transform -1 0 4152 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_187
timestamp 1556798218
transform 1 0 4152 0 1 3810
box 0 0 192 200
use NAND3X1  NAND3X1_2
timestamp 1556798218
transform -1 0 4408 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_70
timestamp 1556798218
transform -1 0 4456 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_113
timestamp 1556798218
transform 1 0 4456 0 1 3810
box 0 0 192 200
use NAND3X1  NAND3X1_3
timestamp 1556798218
transform 1 0 4648 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1556798218
transform -1 0 4776 0 1 3810
box 0 0 64 200
use INVX1  INVX1_7
timestamp 1556798218
transform -1 0 4808 0 1 3810
box 0 0 32 200
use FILL  FILL_19_2_0
timestamp 1556798218
transform 1 0 4808 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1556798218
transform 1 0 4824 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_2
timestamp 1556798218
transform 1 0 4840 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_18
timestamp 1556798218
transform 1 0 4856 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_9
timestamp 1556798218
transform 1 0 4904 0 1 3810
box 0 0 48 200
use INVX1  INVX1_1
timestamp 1556798218
transform -1 0 4984 0 1 3810
box 0 0 32 200
use CLKBUF1  CLKBUF1_25
timestamp 1556798218
transform 1 0 4984 0 1 3810
box 0 0 144 200
use AND2X2  AND2X2_25
timestamp 1556798218
transform 1 0 5128 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_44
timestamp 1556798218
transform -1 0 5256 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_24
timestamp 1556798218
transform -1 0 5304 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_18
timestamp 1556798218
transform 1 0 5304 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_4
timestamp 1556798218
transform -1 0 5432 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_307
timestamp 1556798218
transform 1 0 5432 0 1 3810
box 0 0 192 200
use AND2X2  AND2X2_27
timestamp 1556798218
transform 1 0 5624 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_45
timestamp 1556798218
transform 1 0 5688 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_25
timestamp 1556798218
transform 1 0 5752 0 1 3810
box 0 0 48 200
use INVX1  INVX1_39
timestamp 1556798218
transform -1 0 5832 0 1 3810
box 0 0 32 200
use NAND3X1  NAND3X1_19
timestamp 1556798218
transform 1 0 5832 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1556798218
transform -1 0 5944 0 1 3810
box 0 0 48 200
use OR2X2  OR2X2_5
timestamp 1556798218
transform -1 0 6008 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_161
timestamp 1556798218
transform 1 0 6008 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_478
timestamp 1556798218
transform -1 0 6264 0 1 3810
box 0 0 64 200
use INVX1  INVX1_536
timestamp 1556798218
transform -1 0 6296 0 1 3810
box 0 0 32 200
use FILL  FILL_19_3_0
timestamp 1556798218
transform 1 0 6296 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_1
timestamp 1556798218
transform 1 0 6312 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_2
timestamp 1556798218
transform 1 0 6328 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_315
timestamp 1556798218
transform 1 0 6344 0 1 3810
box 0 0 192 200
use INVX1  INVX1_304
timestamp 1556798218
transform 1 0 6536 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_277
timestamp 1556798218
transform 1 0 6568 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_182
timestamp 1556798218
transform -1 0 6824 0 1 3810
box 0 0 192 200
use BUFX2  BUFX2_6
timestamp 1556798218
transform 1 0 6824 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_279
timestamp 1556798218
transform -1 0 6936 0 1 3810
box 0 0 64 200
use INVX1  INVX1_305
timestamp 1556798218
transform -1 0 6968 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_183
timestamp 1556798218
transform -1 0 7160 0 1 3810
box 0 0 192 200
use CLKBUF1  CLKBUF1_11
timestamp 1556798218
transform -1 0 7304 0 1 3810
box 0 0 144 200
use OAI21X1  OAI21X1_512
timestamp 1556798218
transform 1 0 7304 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_489
timestamp 1556798218
transform -1 0 7416 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_338
timestamp 1556798218
transform 1 0 7416 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_248
timestamp 1556798218
transform -1 0 7656 0 1 3810
box 0 0 48 200
use AND2X2  AND2X2_67
timestamp 1556798218
transform -1 0 7720 0 1 3810
box 0 0 64 200
use INVX1  INVX1_268
timestamp 1556798218
transform 1 0 7720 0 1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_164
timestamp 1556798218
transform -1 0 7944 0 1 3810
box 0 0 192 200
use AOI21X1  AOI21X1_39
timestamp 1556798218
transform -1 0 8008 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_243
timestamp 1556798218
transform -1 0 8072 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_84
timestamp 1556798218
transform 1 0 8072 0 1 3810
box 0 0 64 200
use FILL  FILL_20_1
timestamp 1556798218
transform 1 0 8136 0 1 3810
box 0 0 16 200
use FILL  FILL_20_2
timestamp 1556798218
transform 1 0 8152 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_85
timestamp 1556798218
transform 1 0 8 0 -1 3810
box 0 0 192 200
use INVX1  INVX1_339
timestamp 1556798218
transform 1 0 200 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_308
timestamp 1556798218
transform 1 0 232 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_202
timestamp 1556798218
transform 1 0 296 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_307
timestamp 1556798218
transform -1 0 552 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_338
timestamp 1556798218
transform -1 0 584 0 -1 3810
box 0 0 32 200
use INVX1  INVX1_335
timestamp 1556798218
transform 1 0 584 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_305
timestamp 1556798218
transform -1 0 664 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_306
timestamp 1556798218
transform 1 0 664 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_100
timestamp 1556798218
transform 1 0 712 0 -1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_310
timestamp 1556798218
transform 1 0 792 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_126
timestamp 1556798218
transform -1 0 904 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_101
timestamp 1556798218
transform -1 0 984 0 -1 3810
box 0 0 80 200
use AND2X2  AND2X2_81
timestamp 1556798218
transform -1 0 1048 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_501
timestamp 1556798218
transform -1 0 1096 0 -1 3810
box 0 0 48 200
use AND2X2  AND2X2_134
timestamp 1556798218
transform 1 0 1096 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_232
timestamp 1556798218
transform -1 0 1208 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_231
timestamp 1556798218
transform -1 0 1256 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_61
timestamp 1556798218
transform 1 0 1256 0 -1 3810
box 0 0 192 200
use INVX1  INVX1_83
timestamp 1556798218
transform -1 0 1480 0 -1 3810
box 0 0 32 200
use NOR2X1  NOR2X1_43
timestamp 1556798218
transform -1 0 1528 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_85
timestamp 1556798218
transform 1 0 1528 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_29
timestamp 1556798218
transform -1 0 1672 0 -1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_103
timestamp 1556798218
transform -1 0 1720 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_86
timestamp 1556798218
transform -1 0 1752 0 -1 3810
box 0 0 32 200
use FILL  FILL_18_0_0
timestamp 1556798218
transform 1 0 1752 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1556798218
transform 1 0 1768 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_2
timestamp 1556798218
transform 1 0 1784 0 -1 3810
box 0 0 16 200
use AND2X2  AND2X2_132
timestamp 1556798218
transform 1 0 1800 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_227
timestamp 1556798218
transform -1 0 1912 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_199
timestamp 1556798218
transform 1 0 1912 0 -1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_284
timestamp 1556798218
transform 1 0 2104 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_286
timestamp 1556798218
transform 1 0 2152 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_285
timestamp 1556798218
transform 1 0 2216 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_106
timestamp 1556798218
transform 1 0 2264 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_267
timestamp 1556798218
transform -1 0 2360 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_325
timestamp 1556798218
transform -1 0 2392 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_291
timestamp 1556798218
transform -1 0 2440 0 -1 3810
box 0 0 48 200
use AND2X2  AND2X2_76
timestamp 1556798218
transform 1 0 2440 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_295
timestamp 1556798218
transform 1 0 2504 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_294
timestamp 1556798218
transform -1 0 2600 0 -1 3810
box 0 0 48 200
use BUFX2  BUFX2_18
timestamp 1556798218
transform 1 0 2600 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_316
timestamp 1556798218
transform 1 0 2648 0 -1 3810
box 0 0 32 200
use XNOR2X1  XNOR2X1_42
timestamp 1556798218
transform 1 0 2680 0 -1 3810
box 0 0 112 200
use OAI21X1  OAI21X1_287
timestamp 1556798218
transform 1 0 2792 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_288
timestamp 1556798218
transform -1 0 2920 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_315
timestamp 1556798218
transform 1 0 2920 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_287
timestamp 1556798218
transform -1 0 3000 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_189
timestamp 1556798218
transform 1 0 3000 0 -1 3810
box 0 0 192 200
use INVX1  INVX1_307
timestamp 1556798218
transform 1 0 3192 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_284
timestamp 1556798218
transform -1 0 3288 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_1_0
timestamp 1556798218
transform 1 0 3288 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1556798218
transform 1 0 3304 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_2
timestamp 1556798218
transform 1 0 3320 0 -1 3810
box 0 0 16 200
use NAND3X1  NAND3X1_96
timestamp 1556798218
transform 1 0 3336 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_280
timestamp 1556798218
transform -1 0 3464 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_308
timestamp 1556798218
transform -1 0 3496 0 -1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_45
timestamp 1556798218
transform -1 0 3560 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_500
timestamp 1556798218
transform 1 0 3560 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_279
timestamp 1556798218
transform 1 0 3608 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_283
timestamp 1556798218
transform -1 0 3704 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_310
timestamp 1556798218
transform 1 0 3704 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_188
timestamp 1556798218
transform 1 0 3736 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_328
timestamp 1556798218
transform -1 0 3992 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_361
timestamp 1556798218
transform -1 0 4024 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_215
timestamp 1556798218
transform 1 0 4024 0 -1 3810
box 0 0 192 200
use INVX1  INVX1_355
timestamp 1556798218
transform 1 0 4216 0 -1 3810
box 0 0 32 200
use NOR2X1  NOR2X1_131
timestamp 1556798218
transform -1 0 4296 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_173
timestamp 1556798218
transform 1 0 4296 0 -1 3810
box 0 0 32 200
use AND2X2  AND2X2_18
timestamp 1556798218
transform -1 0 4392 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_585
timestamp 1556798218
transform 1 0 4392 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_343
timestamp 1556798218
transform -1 0 4616 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_520
timestamp 1556798218
transform 1 0 4616 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1556798218
transform -1 0 4728 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_22
timestamp 1556798218
transform 1 0 4728 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_20
timestamp 1556798218
transform -1 0 4824 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_2_0
timestamp 1556798218
transform 1 0 4824 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1556798218
transform 1 0 4840 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_2
timestamp 1556798218
transform 1 0 4856 0 -1 3810
box 0 0 16 200
use NOR2X1  NOR2X1_11
timestamp 1556798218
transform 1 0 4872 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_14
timestamp 1556798218
transform -1 0 4968 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_25
timestamp 1556798218
transform -1 0 5016 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_13
timestamp 1556798218
transform -1 0 5064 0 -1 3810
box 0 0 48 200
use CLKBUF1  CLKBUF1_29
timestamp 1556798218
transform 1 0 5064 0 -1 3810
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_308
timestamp 1556798218
transform 1 0 5208 0 -1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_61
timestamp 1556798218
transform -1 0 5448 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_522
timestamp 1556798218
transform 1 0 5448 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_466
timestamp 1556798218
transform 1 0 5480 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_309
timestamp 1556798218
transform -1 0 5736 0 -1 3810
box 0 0 192 200
use BUFX2  BUFX2_51
timestamp 1556798218
transform 1 0 5736 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_17
timestamp 1556798218
transform -1 0 5832 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_259
timestamp 1556798218
transform 1 0 5832 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_237
timestamp 1556798218
transform -1 0 5928 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_238
timestamp 1556798218
transform -1 0 5992 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_83
timestamp 1556798218
transform -1 0 6056 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_241
timestamp 1556798218
transform 1 0 6056 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_241
timestamp 1556798218
transform -1 0 6168 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_96
timestamp 1556798218
transform 1 0 6168 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_257
timestamp 1556798218
transform -1 0 6248 0 -1 3810
box 0 0 32 200
use AND2X2  AND2X2_73
timestamp 1556798218
transform 1 0 6248 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_277
timestamp 1556798218
transform 1 0 6312 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_3_0
timestamp 1556798218
transform -1 0 6376 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_1
timestamp 1556798218
transform -1 0 6392 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_2
timestamp 1556798218
transform -1 0 6408 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_278
timestamp 1556798218
transform -1 0 6456 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_274
timestamp 1556798218
transform 1 0 6456 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_91
timestamp 1556798218
transform 1 0 6504 0 -1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_110
timestamp 1556798218
transform 1 0 6584 0 -1 3810
box 0 0 48 200
use BUFX2  BUFX2_68
timestamp 1556798218
transform 1 0 6632 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_276
timestamp 1556798218
transform -1 0 6744 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_300
timestamp 1556798218
transform -1 0 6776 0 -1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_276
timestamp 1556798218
transform 1 0 6776 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_90
timestamp 1556798218
transform -1 0 6904 0 -1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_19
timestamp 1556798218
transform -1 0 6952 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_301
timestamp 1556798218
transform -1 0 6984 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_185
timestamp 1556798218
transform -1 0 7176 0 -1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_163
timestamp 1556798218
transform -1 0 7368 0 -1 3810
box 0 0 192 200
use INVX1  INVX1_270
timestamp 1556798218
transform 1 0 7368 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_248
timestamp 1556798218
transform 1 0 7400 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_249
timestamp 1556798218
transform 1 0 7464 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_81
timestamp 1556798218
transform 1 0 7512 0 -1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_99
timestamp 1556798218
transform 1 0 7592 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_245
timestamp 1556798218
transform -1 0 7688 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_269
timestamp 1556798218
transform 1 0 7688 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_246
timestamp 1556798218
transform 1 0 7720 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_245
timestamp 1556798218
transform -1 0 7848 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_80
timestamp 1556798218
transform 1 0 7848 0 -1 3810
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_165
timestamp 1556798218
transform 1 0 7928 0 -1 3810
box 0 0 192 200
use FILL  FILL_19_1
timestamp 1556798218
transform -1 0 8136 0 -1 3810
box 0 0 16 200
use FILL  FILL_19_2
timestamp 1556798218
transform -1 0 8152 0 -1 3810
box 0 0 16 200
use FILL  FILL_19_3
timestamp 1556798218
transform -1 0 8168 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_124
timestamp 1556798218
transform -1 0 72 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_45
timestamp 1556798218
transform 1 0 72 0 1 3410
box 0 0 64 200
use INVX1  INVX1_126
timestamp 1556798218
transform -1 0 168 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_55
timestamp 1556798218
transform 1 0 168 0 1 3410
box 0 0 48 200
use INVX1  INVX1_124
timestamp 1556798218
transform -1 0 248 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_235
timestamp 1556798218
transform 1 0 248 0 1 3410
box 0 0 48 200
use INVX1  INVX1_593
timestamp 1556798218
transform -1 0 328 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_229
timestamp 1556798218
transform -1 0 376 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_230
timestamp 1556798218
transform 1 0 376 0 1 3410
box 0 0 48 200
use AND2X2  AND2X2_133
timestamp 1556798218
transform -1 0 488 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_531
timestamp 1556798218
transform -1 0 552 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_350
timestamp 1556798218
transform 1 0 552 0 1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_203
timestamp 1556798218
transform 1 0 744 0 1 3410
box 0 0 192 200
use INVX1  INVX1_340
timestamp 1556798218
transform -1 0 968 0 1 3410
box 0 0 32 200
use INVX1  INVX1_599
timestamp 1556798218
transform 1 0 968 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_83
timestamp 1556798218
transform 1 0 1000 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_84
timestamp 1556798218
transform -1 0 1128 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_100
timestamp 1556798218
transform -1 0 1176 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_87
timestamp 1556798218
transform 1 0 1176 0 1 3410
box 0 0 64 200
use INVX1  INVX1_84
timestamp 1556798218
transform -1 0 1272 0 1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_33
timestamp 1556798218
transform -1 0 1336 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_32
timestamp 1556798218
transform 1 0 1336 0 1 3410
box 0 0 64 200
use INVX1  INVX1_85
timestamp 1556798218
transform -1 0 1432 0 1 3410
box 0 0 32 200
use AOI22X1  AOI22X1_28
timestamp 1556798218
transform 1 0 1432 0 1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_101
timestamp 1556798218
transform -1 0 1560 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_102
timestamp 1556798218
transform 1 0 1560 0 1 3410
box 0 0 48 200
use AOI21X1  AOI21X1_13
timestamp 1556798218
transform -1 0 1672 0 1 3410
box 0 0 64 200
use XNOR2X1  XNOR2X1_8
timestamp 1556798218
transform -1 0 1784 0 1 3410
box 0 0 112 200
use FILL  FILL_17_0_0
timestamp 1556798218
transform 1 0 1784 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1556798218
transform 1 0 1800 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_2
timestamp 1556798218
transform 1 0 1816 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_60
timestamp 1556798218
transform 1 0 1832 0 1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_191
timestamp 1556798218
transform -1 0 2216 0 1 3410
box 0 0 192 200
use INVX1  INVX1_319
timestamp 1556798218
transform 1 0 2216 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_292
timestamp 1556798218
transform 1 0 2248 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_289
timestamp 1556798218
transform 1 0 2312 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_290
timestamp 1556798218
transform -1 0 2408 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_95
timestamp 1556798218
transform 1 0 2408 0 1 3410
box 0 0 80 200
use NOR2X1  NOR2X1_114
timestamp 1556798218
transform 1 0 2488 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_94
timestamp 1556798218
transform -1 0 2616 0 1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_288
timestamp 1556798218
transform -1 0 2664 0 1 3410
box 0 0 48 200
use INVX1  INVX1_314
timestamp 1556798218
transform 1 0 2664 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_289
timestamp 1556798218
transform 1 0 2696 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_286
timestamp 1556798218
transform 1 0 2760 0 1 3410
box 0 0 48 200
use INVX1  INVX1_306
timestamp 1556798218
transform 1 0 2808 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_111
timestamp 1556798218
transform -1 0 2888 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_281
timestamp 1556798218
transform 1 0 2888 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_97
timestamp 1556798218
transform -1 0 3016 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_280
timestamp 1556798218
transform 1 0 3016 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_216
timestamp 1556798218
transform 1 0 3064 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_319
timestamp 1556798218
transform 1 0 3256 0 1 3410
box 0 0 48 200
use FILL  FILL_17_1_0
timestamp 1556798218
transform 1 0 3304 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1556798218
transform 1 0 3320 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_2
timestamp 1556798218
transform 1 0 3336 0 1 3410
box 0 0 16 200
use INVX1  INVX1_359
timestamp 1556798218
transform 1 0 3352 0 1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_321
timestamp 1556798218
transform 1 0 3384 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_106
timestamp 1556798218
transform -1 0 3512 0 1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_323
timestamp 1556798218
transform 1 0 3512 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_322
timestamp 1556798218
transform 1 0 3560 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_110
timestamp 1556798218
transform -1 0 3672 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_323
timestamp 1556798218
transform 1 0 3672 0 1 3410
box 0 0 64 200
use INVX1  INVX1_357
timestamp 1556798218
transform 1 0 3736 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_324
timestamp 1556798218
transform -1 0 3832 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_111
timestamp 1556798218
transform -1 0 3896 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_217
timestamp 1556798218
transform -1 0 4088 0 1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_342
timestamp 1556798218
transform 1 0 4088 0 1 3410
box 0 0 192 200
use BUFX2  BUFX2_54
timestamp 1556798218
transform 1 0 4280 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_70
timestamp 1556798218
transform -1 0 4376 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_518
timestamp 1556798218
transform -1 0 4440 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_494
timestamp 1556798218
transform -1 0 4488 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_59
timestamp 1556798218
transform 1 0 4488 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_517
timestamp 1556798218
transform -1 0 4616 0 1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_171
timestamp 1556798218
transform -1 0 4696 0 1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_498
timestamp 1556798218
transform 1 0 4696 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_497
timestamp 1556798218
transform -1 0 4792 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_226
timestamp 1556798218
transform 1 0 4792 0 1 3410
box 0 0 48 200
use FILL  FILL_17_2_0
timestamp 1556798218
transform 1 0 4840 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1556798218
transform 1 0 4856 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_2
timestamp 1556798218
transform 1 0 4872 0 1 3410
box 0 0 16 200
use AOI22X1  AOI22X1_170
timestamp 1556798218
transform 1 0 4888 0 1 3410
box 0 0 80 200
use NAND2X1  NAND2X1_496
timestamp 1556798218
transform -1 0 5016 0 1 3410
box 0 0 48 200
use INVX1  INVX1_582
timestamp 1556798218
transform -1 0 5048 0 1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_468
timestamp 1556798218
transform 1 0 5048 0 1 3410
box 0 0 48 200
use XNOR2X1  XNOR2X1_70
timestamp 1556798218
transform 1 0 5096 0 1 3410
box 0 0 112 200
use AOI21X1  AOI21X1_75
timestamp 1556798218
transform 1 0 5208 0 1 3410
box 0 0 64 200
use INVX1  INVX1_519
timestamp 1556798218
transform 1 0 5272 0 1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_156
timestamp 1556798218
transform -1 0 5368 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_449
timestamp 1556798218
transform -1 0 5416 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_152
timestamp 1556798218
transform -1 0 5496 0 1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_461
timestamp 1556798218
transform 1 0 5496 0 1 3410
box 0 0 64 200
use INVX1  INVX1_518
timestamp 1556798218
transform -1 0 5592 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_465
timestamp 1556798218
transform 1 0 5592 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_447
timestamp 1556798218
transform -1 0 5704 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_462
timestamp 1556798218
transform 1 0 5704 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_157
timestamp 1556798218
transform 1 0 5768 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_201
timestamp 1556798218
transform 1 0 5832 0 1 3410
box 0 0 48 200
use INVX1  INVX1_516
timestamp 1556798218
transform -1 0 5912 0 1 3410
box 0 0 32 200
use INVX1  INVX1_260
timestamp 1556798218
transform -1 0 5944 0 1 3410
box 0 0 32 200
use BUFX2  BUFX2_52
timestamp 1556798218
transform 1 0 5944 0 1 3410
box 0 0 48 200
use AND2X2  AND2X2_66
timestamp 1556798218
transform 1 0 5992 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_97
timestamp 1556798218
transform 1 0 6056 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_79
timestamp 1556798218
transform 1 0 6104 0 1 3410
box 0 0 80 200
use AOI22X1  AOI22X1_78
timestamp 1556798218
transform 1 0 6184 0 1 3410
box 0 0 80 200
use NAND3X1  NAND3X1_82
timestamp 1556798218
transform 1 0 6264 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_242
timestamp 1556798218
transform -1 0 6376 0 1 3410
box 0 0 48 200
use FILL  FILL_17_3_0
timestamp 1556798218
transform -1 0 6392 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_1
timestamp 1556798218
transform -1 0 6408 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_2
timestamp 1556798218
transform -1 0 6424 0 1 3410
box 0 0 16 200
use INVX1  INVX1_258
timestamp 1556798218
transform -1 0 6456 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_239
timestamp 1556798218
transform 1 0 6456 0 1 3410
box 0 0 64 200
use INVX1  INVX1_262
timestamp 1556798218
transform 1 0 6520 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_240
timestamp 1556798218
transform 1 0 6552 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_158
timestamp 1556798218
transform -1 0 6808 0 1 3410
box 0 0 192 200
use INVX1  INVX1_302
timestamp 1556798218
transform 1 0 6808 0 1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_94
timestamp 1556798218
transform -1 0 6904 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_274
timestamp 1556798218
transform 1 0 6904 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_275
timestamp 1556798218
transform -1 0 7032 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_275
timestamp 1556798218
transform -1 0 7080 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_278
timestamp 1556798218
transform 1 0 7080 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_95
timestamp 1556798218
transform 1 0 7144 0 1 3410
box 0 0 64 200
use INVX1  INVX1_299
timestamp 1556798218
transform 1 0 7208 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_109
timestamp 1556798218
transform -1 0 7288 0 1 3410
box 0 0 48 200
use INVX1  INVX1_577
timestamp 1556798218
transform 1 0 7288 0 1 3410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_184
timestamp 1556798218
transform -1 0 7512 0 1 3410
box 0 0 192 200
use CLKBUF1  CLKBUF1_38
timestamp 1556798218
transform -1 0 7656 0 1 3410
box 0 0 144 200
use INVX1  INVX1_273
timestamp 1556798218
transform 1 0 7656 0 1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_255
timestamp 1556798218
transform 1 0 7688 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_256
timestamp 1556798218
transform -1 0 7784 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_162
timestamp 1556798218
transform -1 0 7976 0 1 3410
box 0 0 192 200
use CLKBUF1  CLKBUF1_46
timestamp 1556798218
transform 1 0 7976 0 1 3410
box 0 0 144 200
use FILL  FILL_18_1
timestamp 1556798218
transform 1 0 8120 0 1 3410
box 0 0 16 200
use FILL  FILL_18_2
timestamp 1556798218
transform 1 0 8136 0 1 3410
box 0 0 16 200
use FILL  FILL_18_3
timestamp 1556798218
transform 1 0 8152 0 1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_19
timestamp 1556798218
transform -1 0 72 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_44
timestamp 1556798218
transform 1 0 72 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_134
timestamp 1556798218
transform -1 0 184 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_121
timestamp 1556798218
transform 1 0 184 0 -1 3410
box 0 0 64 200
use XNOR2X1  XNOR2X1_14
timestamp 1556798218
transform -1 0 360 0 -1 3410
box 0 0 112 200
use INVX1  INVX1_127
timestamp 1556798218
transform 1 0 360 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_120
timestamp 1556798218
transform -1 0 456 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_508
timestamp 1556798218
transform 1 0 456 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_179
timestamp 1556798218
transform 1 0 504 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_528
timestamp 1556798218
transform 1 0 568 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_527
timestamp 1556798218
transform -1 0 696 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_595
timestamp 1556798218
transform -1 0 728 0 -1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_178
timestamp 1556798218
transform 1 0 728 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_529
timestamp 1556798218
transform -1 0 856 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_594
timestamp 1556798218
transform -1 0 888 0 -1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_509
timestamp 1556798218
transform 1 0 888 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_174
timestamp 1556798218
transform -1 0 1016 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_532
timestamp 1556798218
transform 1 0 1016 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_351
timestamp 1556798218
transform 1 0 1080 0 -1 3410
box 0 0 192 200
use BUFX2  BUFX2_117
timestamp 1556798218
transform -1 0 1320 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_341
timestamp 1556798218
transform 1 0 1320 0 -1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_127
timestamp 1556798218
transform -1 0 1400 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_209
timestamp 1556798218
transform -1 0 1592 0 -1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_107
timestamp 1556798218
transform 1 0 1592 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_312
timestamp 1556798218
transform -1 0 1720 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_42
timestamp 1556798218
transform -1 0 1768 0 -1 3410
box 0 0 48 200
use FILL  FILL_16_0_0
timestamp 1556798218
transform -1 0 1784 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1556798218
transform -1 0 1800 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_2
timestamp 1556798218
transform -1 0 1816 0 -1 3410
box 0 0 16 200
use INVX1  INVX1_82
timestamp 1556798218
transform -1 0 1848 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_88
timestamp 1556798218
transform -1 0 1912 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_88
timestamp 1556798218
transform -1 0 1944 0 -1 3410
box 0 0 32 200
use BUFX2  BUFX2_76
timestamp 1556798218
transform -1 0 1992 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_59
timestamp 1556798218
transform 1 0 1992 0 -1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_325
timestamp 1556798218
transform 1 0 2184 0 -1 3410
box 0 0 192 200
use BUFX2  BUFX2_74
timestamp 1556798218
transform 1 0 2376 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_165
timestamp 1556798218
transform -1 0 2488 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_486
timestamp 1556798218
transform -1 0 2552 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_485
timestamp 1556798218
transform 1 0 2552 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_546
timestamp 1556798218
transform 1 0 2616 0 -1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_470
timestamp 1556798218
transform -1 0 2696 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_489
timestamp 1556798218
transform 1 0 2696 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_544
timestamp 1556798218
transform -1 0 2792 0 -1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_215
timestamp 1556798218
transform -1 0 2840 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_290
timestamp 1556798218
transform -1 0 2904 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_318
timestamp 1556798218
transform -1 0 2936 0 -1 3410
box 0 0 32 200
use AND2X2  AND2X2_75
timestamp 1556798218
transform -1 0 3000 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_190
timestamp 1556798218
transform -1 0 3192 0 -1 3410
box 0 0 192 200
use AND2X2  AND2X2_12
timestamp 1556798218
transform -1 0 3256 0 -1 3410
box 0 0 64 200
use BUFX2  BUFX2_122
timestamp 1556798218
transform 1 0 3256 0 -1 3410
box 0 0 48 200
use FILL  FILL_16_1_0
timestamp 1556798218
transform 1 0 3304 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1556798218
transform 1 0 3320 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_2
timestamp 1556798218
transform 1 0 3336 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_84
timestamp 1556798218
transform 1 0 3352 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_360
timestamp 1556798218
transform 1 0 3416 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_326
timestamp 1556798218
transform 1 0 3448 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_214
timestamp 1556798218
transform 1 0 3512 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_325
timestamp 1556798218
transform -1 0 3768 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_107
timestamp 1556798218
transform 1 0 3768 0 -1 3410
box 0 0 80 200
use INVX1  INVX1_358
timestamp 1556798218
transform 1 0 3848 0 -1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_132
timestamp 1556798218
transform -1 0 3928 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_356
timestamp 1556798218
transform 1 0 3928 0 -1 3410
box 0 0 32 200
use AOI21X1  AOI21X1_52
timestamp 1556798218
transform 1 0 3960 0 -1 3410
box 0 0 64 200
use XNOR2X1  XNOR2X1_47
timestamp 1556798218
transform -1 0 4136 0 -1 3410
box 0 0 112 200
use OAI21X1  OAI21X1_327
timestamp 1556798218
transform 1 0 4136 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_320
timestamp 1556798218
transform -1 0 4248 0 -1 3410
box 0 0 48 200
use BUFX2  BUFX2_127
timestamp 1556798218
transform -1 0 4296 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_178
timestamp 1556798218
transform 1 0 4296 0 -1 3410
box 0 0 32 200
use AND2X2  AND2X2_52
timestamp 1556798218
transform 1 0 4328 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_344
timestamp 1556798218
transform -1 0 4584 0 -1 3410
box 0 0 192 200
use INVX1  INVX1_583
timestamp 1556798218
transform 1 0 4584 0 -1 3410
box 0 0 32 200
use XNOR2X1  XNOR2X1_79
timestamp 1556798218
transform 1 0 4616 0 -1 3410
box 0 0 112 200
use AOI21X1  AOI21X1_84
timestamp 1556798218
transform 1 0 4728 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_584
timestamp 1556798218
transform -1 0 4824 0 -1 3410
box 0 0 32 200
use FILL  FILL_16_2_0
timestamp 1556798218
transform -1 0 4840 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1556798218
transform -1 0 4856 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_2
timestamp 1556798218
transform -1 0 4872 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_131
timestamp 1556798218
transform -1 0 4936 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_580
timestamp 1556798218
transform 1 0 4936 0 -1 3410
box 0 0 32 200
use BUFX2  BUFX2_128
timestamp 1556798218
transform 1 0 4968 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_174
timestamp 1556798218
transform 1 0 5016 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_516
timestamp 1556798218
transform 1 0 5080 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_495
timestamp 1556798218
transform 1 0 5144 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_519
timestamp 1556798218
transform -1 0 5256 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_581
timestamp 1556798218
transform 1 0 5256 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_515
timestamp 1556798218
transform -1 0 5352 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_450
timestamp 1556798218
transform 1 0 5352 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_448
timestamp 1556798218
transform 1 0 5400 0 -1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_202
timestamp 1556798218
transform 1 0 5448 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_153
timestamp 1556798218
transform 1 0 5496 0 -1 3410
box 0 0 80 200
use INVX1  INVX1_520
timestamp 1556798218
transform 1 0 5576 0 -1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_446
timestamp 1556798218
transform -1 0 5656 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_517
timestamp 1556798218
transform 1 0 5656 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_463
timestamp 1556798218
transform 1 0 5688 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_464
timestamp 1556798218
transform -1 0 5816 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_306
timestamp 1556798218
transform -1 0 6008 0 -1 3410
box 0 0 192 200
use AND2X2  AND2X2_130
timestamp 1556798218
transform 1 0 6008 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_243
timestamp 1556798218
transform 1 0 6072 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_244
timestamp 1556798218
transform -1 0 6168 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_160
timestamp 1556798218
transform -1 0 6360 0 -1 3410
box 0 0 192 200
use FILL  FILL_16_3_0
timestamp 1556798218
transform -1 0 6376 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_1
timestamp 1556798218
transform -1 0 6392 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_2
timestamp 1556798218
transform -1 0 6408 0 -1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_38
timestamp 1556798218
transform -1 0 6472 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_261
timestamp 1556798218
transform -1 0 6504 0 -1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_240
timestamp 1556798218
transform -1 0 6552 0 -1 3410
box 0 0 48 200
use XNOR2X1  XNOR2X1_33
timestamp 1556798218
transform 1 0 6552 0 -1 3410
box 0 0 112 200
use AND2X2  AND2X2_71
timestamp 1556798218
transform -1 0 6728 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_303
timestamp 1556798218
transform -1 0 6760 0 -1 3410
box 0 0 32 200
use CLKBUF1  CLKBUF1_37
timestamp 1556798218
transform -1 0 6904 0 -1 3410
box 0 0 144 200
use XNOR2X1  XNOR2X1_39
timestamp 1556798218
transform -1 0 7016 0 -1 3410
box 0 0 112 200
use AOI21X1  AOI21X1_44
timestamp 1556798218
transform 1 0 7016 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_292
timestamp 1556798218
transform 1 0 7080 0 -1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_107
timestamp 1556798218
transform -1 0 7160 0 -1 3410
box 0 0 48 200
use BUFX2  BUFX2_124
timestamp 1556798218
transform 1 0 7160 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_271
timestamp 1556798218
transform 1 0 7208 0 -1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_100
timestamp 1556798218
transform -1 0 7288 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_169
timestamp 1556798218
transform -1 0 7480 0 -1 3410
box 0 0 192 200
use INVX1  INVX1_33
timestamp 1556798218
transform -1 0 7512 0 -1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_87
timestamp 1556798218
transform 1 0 7512 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_274
timestamp 1556798218
transform -1 0 7608 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_251
timestamp 1556798218
transform 1 0 7608 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_250
timestamp 1556798218
transform 1 0 7672 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_254
timestamp 1556798218
transform -1 0 7800 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_253
timestamp 1556798218
transform -1 0 7848 0 -1 3410
box 0 0 48 200
use XNOR2X1  XNOR2X1_35
timestamp 1556798218
transform -1 0 7960 0 -1 3410
box 0 0 112 200
use AOI21X1  AOI21X1_40
timestamp 1556798218
transform -1 0 8024 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_275
timestamp 1556798218
transform -1 0 8056 0 -1 3410
box 0 0 32 200
use BUFX2  BUFX2_138
timestamp 1556798218
transform 1 0 8056 0 -1 3410
box 0 0 48 200
use BUFX2  BUFX2_140
timestamp 1556798218
transform 1 0 8104 0 -1 3410
box 0 0 48 200
use FILL  FILL_17_1
timestamp 1556798218
transform -1 0 8168 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_135
timestamp 1556798218
transform 1 0 8 0 1 3010
box 0 0 48 200
use INVX1  INVX1_125
timestamp 1556798218
transform 1 0 56 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_40
timestamp 1556798218
transform -1 0 168 0 1 3010
box 0 0 80 200
use AND2X2  AND2X2_44
timestamp 1556798218
transform 1 0 168 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_56
timestamp 1556798218
transform -1 0 280 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_136
timestamp 1556798218
transform 1 0 280 0 1 3010
box 0 0 48 200
use BUFX2  BUFX2_82
timestamp 1556798218
transform -1 0 376 0 1 3010
box 0 0 48 200
use BUFX2  BUFX2_78
timestamp 1556798218
transform 1 0 376 0 1 3010
box 0 0 48 200
use XNOR2X1  XNOR2X1_81
timestamp 1556798218
transform 1 0 424 0 1 3010
box 0 0 112 200
use AOI21X1  AOI21X1_86
timestamp 1556798218
transform -1 0 600 0 1 3010
box 0 0 64 200
use INVX1  INVX1_597
timestamp 1556798218
transform -1 0 632 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_507
timestamp 1556798218
transform -1 0 680 0 1 3010
box 0 0 48 200
use INVX1  INVX1_596
timestamp 1556798218
transform 1 0 680 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_530
timestamp 1556798218
transform 1 0 712 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_236
timestamp 1556798218
transform -1 0 824 0 1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_175
timestamp 1556798218
transform -1 0 904 0 1 3010
box 0 0 80 200
use CLKBUF1  CLKBUF1_14
timestamp 1556798218
transform 1 0 904 0 1 3010
box 0 0 144 200
use XNOR2X1  XNOR2X1_45
timestamp 1556798218
transform 1 0 1048 0 1 3010
box 0 0 112 200
use AOI21X1  AOI21X1_50
timestamp 1556798218
transform 1 0 1160 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_301
timestamp 1556798218
transform -1 0 1272 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_315
timestamp 1556798218
transform -1 0 1336 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_310
timestamp 1556798218
transform -1 0 1384 0 1 3010
box 0 0 48 200
use INVX1  INVX1_342
timestamp 1556798218
transform 1 0 1384 0 1 3010
box 0 0 32 200
use INVX1  INVX1_343
timestamp 1556798218
transform -1 0 1448 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_311
timestamp 1556798218
transform -1 0 1512 0 1 3010
box 0 0 64 200
use INVX1  INVX1_344
timestamp 1556798218
transform 1 0 1512 0 1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_106
timestamp 1556798218
transform -1 0 1608 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_311
timestamp 1556798218
transform 1 0 1608 0 1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_102
timestamp 1556798218
transform -1 0 1736 0 1 3010
box 0 0 80 200
use FILL  FILL_15_0_0
timestamp 1556798218
transform -1 0 1752 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1556798218
transform -1 0 1768 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_2
timestamp 1556798218
transform -1 0 1784 0 1 3010
box 0 0 16 200
use NOR2X1  NOR2X1_128
timestamp 1556798218
transform -1 0 1832 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_313
timestamp 1556798218
transform 1 0 1832 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_312
timestamp 1556798218
transform -1 0 1928 0 1 3010
box 0 0 48 200
use BUFX2  BUFX2_77
timestamp 1556798218
transform -1 0 1976 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_3
timestamp 1556798218
transform 1 0 1976 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_2
timestamp 1556798218
transform 1 0 2024 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_4
timestamp 1556798218
transform -1 0 2120 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_322
timestamp 1556798218
transform 1 0 2120 0 1 3010
box 0 0 192 200
use INVX1  INVX1_549
timestamp 1556798218
transform 1 0 2312 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_488
timestamp 1556798218
transform 1 0 2344 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_487
timestamp 1556798218
transform -1 0 2472 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_164
timestamp 1556798218
transform 1 0 2472 0 1 3010
box 0 0 64 200
use INVX1  INVX1_545
timestamp 1556798218
transform -1 0 2568 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_160
timestamp 1556798218
transform -1 0 2648 0 1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_471
timestamp 1556798218
transform -1 0 2696 0 1 3010
box 0 0 48 200
use INVX1  INVX1_548
timestamp 1556798218
transform 1 0 2696 0 1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_79
timestamp 1556798218
transform -1 0 2792 0 1 3010
box 0 0 64 200
use XNOR2X1  XNOR2X1_74
timestamp 1556798218
transform -1 0 2904 0 1 3010
box 0 0 112 200
use INVX1  INVX1_606
timestamp 1556798218
transform 1 0 2904 0 1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_355
timestamp 1556798218
transform -1 0 3128 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_538
timestamp 1556798218
transform 1 0 3128 0 1 3010
box 0 0 64 200
use FILL  FILL_15_1_0
timestamp 1556798218
transform 1 0 3192 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1556798218
transform 1 0 3208 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_2
timestamp 1556798218
transform 1 0 3224 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_354
timestamp 1556798218
transform 1 0 3240 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_536
timestamp 1556798218
transform 1 0 3432 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_535
timestamp 1556798218
transform -1 0 3560 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_177
timestamp 1556798218
transform -1 0 3640 0 1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_512
timestamp 1556798218
transform -1 0 3688 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_516
timestamp 1556798218
transform 1 0 3688 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_515
timestamp 1556798218
transform -1 0 3784 0 1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_87
timestamp 1556798218
transform 1 0 3784 0 1 3010
box 0 0 64 200
use INVX1  INVX1_604
timestamp 1556798218
transform 1 0 3848 0 1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_356
timestamp 1556798218
transform -1 0 4072 0 1 3010
box 0 0 192 200
use CLKBUF1  CLKBUF1_32
timestamp 1556798218
transform -1 0 4216 0 1 3010
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_112
timestamp 1556798218
transform 1 0 4216 0 1 3010
box 0 0 192 200
use INVX1  INVX1_174
timestamp 1556798218
transform 1 0 4408 0 1 3010
box 0 0 32 200
use INVX1  INVX1_175
timestamp 1556798218
transform 1 0 4440 0 1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_58
timestamp 1556798218
transform -1 0 4536 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_164
timestamp 1556798218
transform 1 0 4536 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_163
timestamp 1556798218
transform -1 0 4664 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_173
timestamp 1556798218
transform -1 0 4712 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_167
timestamp 1556798218
transform 1 0 4712 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_213
timestamp 1556798218
transform 1 0 4776 0 1 3010
box 0 0 48 200
use FILL  FILL_15_2_0
timestamp 1556798218
transform 1 0 4824 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1556798218
transform 1 0 4840 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_2
timestamp 1556798218
transform 1 0 4856 0 1 3010
box 0 0 16 200
use NOR2X1  NOR2X1_214
timestamp 1556798218
transform 1 0 4872 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_211
timestamp 1556798218
transform 1 0 4920 0 1 3010
box 0 0 48 200
use AND2X2  AND2X2_124
timestamp 1556798218
transform 1 0 4968 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_212
timestamp 1556798218
transform -1 0 5080 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_175
timestamp 1556798218
transform -1 0 5144 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_345
timestamp 1556798218
transform 1 0 5144 0 1 3010
box 0 0 192 200
use NOR2X1  NOR2X1_225
timestamp 1556798218
transform 1 0 5336 0 1 3010
box 0 0 48 200
use INVX1  INVX1_579
timestamp 1556798218
transform -1 0 5416 0 1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_217
timestamp 1556798218
transform 1 0 5416 0 1 3010
box 0 0 48 200
use INVX1  INVX1_551
timestamp 1556798218
transform -1 0 5496 0 1 3010
box 0 0 32 200
use AND2X2  AND2X2_119
timestamp 1556798218
transform -1 0 5560 0 1 3010
box 0 0 64 200
use XNOR2X1  XNOR2X1_75
timestamp 1556798218
transform -1 0 5672 0 1 3010
box 0 0 112 200
use BUFX2  BUFX2_93
timestamp 1556798218
transform -1 0 5720 0 1 3010
box 0 0 48 200
use BUFX2  BUFX2_94
timestamp 1556798218
transform -1 0 5768 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_12
timestamp 1556798218
transform -1 0 5816 0 1 3010
box 0 0 48 200
use INVX1  INVX1_521
timestamp 1556798218
transform -1 0 5848 0 1 3010
box 0 0 32 200
use BUFX2  BUFX2_33
timestamp 1556798218
transform -1 0 5896 0 1 3010
box 0 0 48 200
use BUFX2  BUFX2_126
timestamp 1556798218
transform -1 0 5944 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_159
timestamp 1556798218
transform -1 0 6136 0 1 3010
box 0 0 192 200
use INVX1  INVX1_263
timestamp 1556798218
transform 1 0 6136 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_242
timestamp 1556798218
transform -1 0 6232 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_64
timestamp 1556798218
transform -1 0 6296 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_273
timestamp 1556798218
transform 1 0 6296 0 1 3010
box 0 0 48 200
use FILL  FILL_15_3_0
timestamp 1556798218
transform -1 0 6360 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_1
timestamp 1556798218
transform -1 0 6376 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_2
timestamp 1556798218
transform -1 0 6392 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_272
timestamp 1556798218
transform -1 0 6440 0 1 3010
box 0 0 48 200
use AND2X2  AND2X2_72
timestamp 1556798218
transform 1 0 6440 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_89
timestamp 1556798218
transform 1 0 6504 0 1 3010
box 0 0 80 200
use NOR2X1  NOR2X1_108
timestamp 1556798218
transform 1 0 6584 0 1 3010
box 0 0 48 200
use INVX1  INVX1_295
timestamp 1556798218
transform 1 0 6632 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_88
timestamp 1556798218
transform -1 0 6744 0 1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_271
timestamp 1556798218
transform 1 0 6744 0 1 3010
box 0 0 48 200
use INVX1  INVX1_297
timestamp 1556798218
transform 1 0 6792 0 1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_92
timestamp 1556798218
transform -1 0 6888 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_268
timestamp 1556798218
transform 1 0 6888 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_269
timestamp 1556798218
transform -1 0 7016 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_93
timestamp 1556798218
transform -1 0 7080 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_272
timestamp 1556798218
transform -1 0 7144 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_270
timestamp 1556798218
transform -1 0 7192 0 1 3010
box 0 0 48 200
use INVX1  INVX1_294
timestamp 1556798218
transform -1 0 7224 0 1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_181
timestamp 1556798218
transform -1 0 7416 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_254
timestamp 1556798218
transform 1 0 7416 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_86
timestamp 1556798218
transform -1 0 7528 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_82
timestamp 1556798218
transform -1 0 7608 0 1 3010
box 0 0 80 200
use NOR2X1  NOR2X1_101
timestamp 1556798218
transform -1 0 7656 0 1 3010
box 0 0 48 200
use INVX1  INVX1_272
timestamp 1556798218
transform -1 0 7688 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_252
timestamp 1556798218
transform 1 0 7688 0 1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_83
timestamp 1556798218
transform 1 0 7736 0 1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_252
timestamp 1556798218
transform 1 0 7816 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_255
timestamp 1556798218
transform 1 0 7880 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_167
timestamp 1556798218
transform -1 0 8136 0 1 3010
box 0 0 192 200
use FILL  FILL_16_1
timestamp 1556798218
transform 1 0 8136 0 1 3010
box 0 0 16 200
use FILL  FILL_16_2
timestamp 1556798218
transform 1 0 8152 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_133
timestamp 1556798218
transform 1 0 8 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_128
timestamp 1556798218
transform -1 0 88 0 -1 3010
box 0 0 32 200
use INVX1  INVX1_129
timestamp 1556798218
transform 1 0 88 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_123
timestamp 1556798218
transform 1 0 120 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_122
timestamp 1556798218
transform 1 0 184 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_41
timestamp 1556798218
transform -1 0 328 0 -1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_137
timestamp 1556798218
transform -1 0 376 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_352
timestamp 1556798218
transform 1 0 376 0 -1 3010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_353
timestamp 1556798218
transform 1 0 568 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_598
timestamp 1556798218
transform -1 0 792 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_511
timestamp 1556798218
transform 1 0 792 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_510
timestamp 1556798218
transform -1 0 888 0 -1 3010
box 0 0 48 200
use AND2X2  AND2X2_136
timestamp 1556798218
transform -1 0 952 0 -1 3010
box 0 0 64 200
use CLKBUF1  CLKBUF1_41
timestamp 1556798218
transform 1 0 952 0 -1 3010
box 0 0 144 200
use BUFX2  BUFX2_81
timestamp 1556798218
transform -1 0 1144 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_208
timestamp 1556798218
transform 1 0 1144 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_345
timestamp 1556798218
transform 1 0 1336 0 -1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_206
timestamp 1556798218
transform 1 0 1368 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_313
timestamp 1556798218
transform 1 0 1560 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_314
timestamp 1556798218
transform -1 0 1688 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_346
timestamp 1556798218
transform -1 0 1720 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_309
timestamp 1556798218
transform -1 0 1768 0 -1 3010
box 0 0 48 200
use FILL  FILL_14_0_0
timestamp 1556798218
transform -1 0 1784 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1556798218
transform -1 0 1800 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_2
timestamp 1556798218
transform -1 0 1816 0 -1 3010
box 0 0 16 200
use AOI22X1  AOI22X1_103
timestamp 1556798218
transform -1 0 1896 0 -1 3010
box 0 0 80 200
use AND2X2  AND2X2_82
timestamp 1556798218
transform -1 0 1960 0 -1 3010
box 0 0 64 200
use BUFX2  BUFX2_73
timestamp 1556798218
transform -1 0 2008 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_316
timestamp 1556798218
transform -1 0 2072 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_347
timestamp 1556798218
transform -1 0 2104 0 -1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_207
timestamp 1556798218
transform 1 0 2104 0 -1 3010
box 0 0 192 200
use BUFX2  BUFX2_75
timestamp 1556798218
transform -1 0 2344 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_469
timestamp 1556798218
transform 1 0 2344 0 -1 3010
box 0 0 48 200
use AND2X2  AND2X2_126
timestamp 1556798218
transform 1 0 2392 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_216
timestamp 1556798218
transform -1 0 2504 0 -1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_161
timestamp 1556798218
transform -1 0 2584 0 -1 3010
box 0 0 80 200
use INVX1  INVX1_547
timestamp 1556798218
transform -1 0 2616 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_472
timestamp 1556798218
transform 1 0 2616 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_473
timestamp 1556798218
transform -1 0 2712 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_324
timestamp 1556798218
transform 1 0 2712 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_490
timestamp 1556798218
transform -1 0 2968 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_550
timestamp 1556798218
transform -1 0 3000 0 -1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_323
timestamp 1556798218
transform 1 0 3000 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_600
timestamp 1556798218
transform 1 0 3192 0 -1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_237
timestamp 1556798218
transform -1 0 3272 0 -1 3010
box 0 0 48 200
use FILL  FILL_14_1_0
timestamp 1556798218
transform 1 0 3272 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1556798218
transform 1 0 3288 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_2
timestamp 1556798218
transform 1 0 3304 0 -1 3010
box 0 0 16 200
use AOI22X1  AOI22X1_176
timestamp 1556798218
transform 1 0 3320 0 -1 3010
box 0 0 80 200
use INVX1  INVX1_603
timestamp 1556798218
transform 1 0 3400 0 -1 3010
box 0 0 32 200
use INVX1  INVX1_605
timestamp 1556798218
transform -1 0 3464 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_514
timestamp 1556798218
transform -1 0 3512 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_601
timestamp 1556798218
transform -1 0 3544 0 -1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_238
timestamp 1556798218
transform 1 0 3544 0 -1 3010
box 0 0 48 200
use AND2X2  AND2X2_137
timestamp 1556798218
transform -1 0 3656 0 -1 3010
box 0 0 64 200
use XNOR2X1  XNOR2X1_82
timestamp 1556798218
transform 1 0 3656 0 -1 3010
box 0 0 112 200
use NAND2X1  NAND2X1_513
timestamp 1556798218
transform 1 0 3768 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_537
timestamp 1556798218
transform -1 0 3880 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_602
timestamp 1556798218
transform 1 0 3880 0 -1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_181
timestamp 1556798218
transform 1 0 3912 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_534
timestamp 1556798218
transform 1 0 3976 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_533
timestamp 1556798218
transform -1 0 4104 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_180
timestamp 1556798218
transform 1 0 4104 0 -1 3010
box 0 0 64 200
use BUFX2  BUFX2_102
timestamp 1556798218
transform -1 0 4216 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_110
timestamp 1556798218
transform 1 0 4216 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_166
timestamp 1556798218
transform 1 0 4408 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_165
timestamp 1556798218
transform -1 0 4536 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_172
timestamp 1556798218
transform -1 0 4584 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_177
timestamp 1556798218
transform 1 0 4584 0 -1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_54
timestamp 1556798218
transform 1 0 4616 0 -1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_174
timestamp 1556798218
transform -1 0 4744 0 -1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_26
timestamp 1556798218
transform -1 0 4808 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_2_0
timestamp 1556798218
transform -1 0 4824 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1556798218
transform -1 0 4840 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_2
timestamp 1556798218
transform -1 0 4856 0 -1 3010
box 0 0 16 200
use XNOR2X1  XNOR2X1_21
timestamp 1556798218
transform -1 0 4968 0 -1 3010
box 0 0 112 200
use AND2X2  AND2X2_125
timestamp 1556798218
transform -1 0 5032 0 -1 3010
box 0 0 64 200
use BUFX2  BUFX2_99
timestamp 1556798218
transform -1 0 5080 0 -1 3010
box 0 0 48 200
use NOR3X1  NOR3X1_7
timestamp 1556798218
transform -1 0 5208 0 -1 3010
box 0 0 128 200
use NAND2X1  NAND2X1_466
timestamp 1556798218
transform -1 0 5256 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_555
timestamp 1556798218
transform 1 0 5256 0 -1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_328
timestamp 1556798218
transform 1 0 5288 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_554
timestamp 1556798218
transform 1 0 5480 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_80
timestamp 1556798218
transform 1 0 5512 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_495
timestamp 1556798218
transform -1 0 5640 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_553
timestamp 1556798218
transform -1 0 5672 0 -1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_166
timestamp 1556798218
transform -1 0 5736 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_167
timestamp 1556798218
transform 1 0 5736 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_329
timestamp 1556798218
transform -1 0 5992 0 -1 3010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_155
timestamp 1556798218
transform -1 0 6184 0 -1 3010
box 0 0 192 200
use AND2X2  AND2X2_14
timestamp 1556798218
transform 1 0 6184 0 -1 3010
box 0 0 64 200
use BUFX2  BUFX2_100
timestamp 1556798218
transform 1 0 6248 0 -1 3010
box 0 0 48 200
use FILL  FILL_14_3_0
timestamp 1556798218
transform -1 0 6312 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_1
timestamp 1556798218
transform -1 0 6328 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_2
timestamp 1556798218
transform -1 0 6344 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_179
timestamp 1556798218
transform -1 0 6536 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_298
timestamp 1556798218
transform 1 0 6536 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_273
timestamp 1556798218
transform -1 0 6632 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_178
timestamp 1556798218
transform -1 0 6824 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_271
timestamp 1556798218
transform 1 0 6824 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_270
timestamp 1556798218
transform -1 0 6952 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_269
timestamp 1556798218
transform -1 0 7000 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_296
timestamp 1556798218
transform 1 0 7000 0 -1 3010
box 0 0 32 200
use INVX1  INVX1_293
timestamp 1556798218
transform 1 0 7032 0 -1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_43
timestamp 1556798218
transform 1 0 7064 0 -1 3010
box 0 0 64 200
use XNOR2X1  XNOR2X1_38
timestamp 1556798218
transform -1 0 7240 0 -1 3010
box 0 0 112 200
use CLKBUF1  CLKBUF1_20
timestamp 1556798218
transform -1 0 7384 0 -1 3010
box 0 0 144 200
use NAND2X1  NAND2X1_45
timestamp 1556798218
transform 1 0 7384 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_28
timestamp 1556798218
transform 1 0 7432 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1556798218
transform -1 0 7528 0 -1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1556798218
transform -1 0 7720 0 -1 3010
box 0 0 192 200
use AND2X2  AND2X2_68
timestamp 1556798218
transform 1 0 7720 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_276
timestamp 1556798218
transform 1 0 7784 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_253
timestamp 1556798218
transform 1 0 7816 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_166
timestamp 1556798218
transform 1 0 7880 0 -1 3010
box 0 0 192 200
use BUFX2  BUFX2_143
timestamp 1556798218
transform 1 0 8072 0 -1 3010
box 0 0 48 200
use FILL  FILL_15_1
timestamp 1556798218
transform -1 0 8136 0 -1 3010
box 0 0 16 200
use FILL  FILL_15_2
timestamp 1556798218
transform -1 0 8152 0 -1 3010
box 0 0 16 200
use FILL  FILL_15_3
timestamp 1556798218
transform -1 0 8168 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_84
timestamp 1556798218
transform 1 0 8 0 1 2610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_82
timestamp 1556798218
transform -1 0 392 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_125
timestamp 1556798218
transform -1 0 456 0 1 2610
box 0 0 64 200
use INVX1  INVX1_130
timestamp 1556798218
transform -1 0 488 0 1 2610
box 0 0 32 200
use AND2X2  AND2X2_139
timestamp 1556798218
transform 1 0 488 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_83
timestamp 1556798218
transform 1 0 552 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_5
timestamp 1556798218
transform -1 0 792 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_3
timestamp 1556798218
transform 1 0 792 0 1 2610
box 0 0 48 200
use BUFX2  BUFX2_13
timestamp 1556798218
transform -1 0 888 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_6
timestamp 1556798218
transform -1 0 936 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_145
timestamp 1556798218
transform 1 0 936 0 1 2610
box 0 0 48 200
use INVX1  INVX1_383
timestamp 1556798218
transform -1 0 1016 0 1 2610
box 0 0 32 200
use AOI21X1  AOI21X1_56
timestamp 1556798218
transform -1 0 1080 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_344
timestamp 1556798218
transform 1 0 1080 0 1 2610
box 0 0 48 200
use XNOR2X1  XNOR2X1_51
timestamp 1556798218
transform -1 0 1240 0 1 2610
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_226
timestamp 1556798218
transform 1 0 1240 0 1 2610
box 0 0 192 200
use CLKBUF1  CLKBUF1_48
timestamp 1556798218
transform 1 0 1432 0 1 2610
box 0 0 144 200
use OAI21X1  OAI21X1_343
timestamp 1556798218
transform -1 0 1640 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_344
timestamp 1556798218
transform -1 0 1704 0 1 2610
box 0 0 64 200
use INVX1  INVX1_381
timestamp 1556798218
transform -1 0 1736 0 1 2610
box 0 0 32 200
use FILL  FILL_13_0_0
timestamp 1556798218
transform -1 0 1752 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1556798218
transform -1 0 1768 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_2
timestamp 1556798218
transform -1 0 1784 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_337
timestamp 1556798218
transform -1 0 1832 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_339
timestamp 1556798218
transform 1 0 1832 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_90
timestamp 1556798218
transform -1 0 1944 0 1 2610
box 0 0 64 200
use INVX1  INVX1_377
timestamp 1556798218
transform 1 0 1944 0 1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_338
timestamp 1556798218
transform -1 0 2024 0 1 2610
box 0 0 48 200
use AOI21X1  AOI21X1_55
timestamp 1556798218
transform -1 0 2088 0 1 2610
box 0 0 64 200
use BUFX2  BUFX2_36
timestamp 1556798218
transform 1 0 2088 0 1 2610
box 0 0 48 200
use XNOR2X1  XNOR2X1_50
timestamp 1556798218
transform -1 0 2248 0 1 2610
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_228
timestamp 1556798218
transform -1 0 2440 0 1 2610
box 0 0 192 200
use BUFX2  BUFX2_3
timestamp 1556798218
transform -1 0 2488 0 1 2610
box 0 0 48 200
use CLKBUF1  CLKBUF1_19
timestamp 1556798218
transform 1 0 2488 0 1 2610
box 0 0 144 200
use NOR2X1  NOR2X1_120
timestamp 1556798218
transform 1 0 2632 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_67
timestamp 1556798218
transform 1 0 2680 0 1 2610
box 0 0 192 200
use BUFX2  BUFX2_27
timestamp 1556798218
transform -1 0 2920 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_295
timestamp 1556798218
transform -1 0 3112 0 1 2610
box 0 0 192 200
use INVX1  INVX1_501
timestamp 1556798218
transform 1 0 3112 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_448
timestamp 1556798218
transform 1 0 3144 0 1 2610
box 0 0 64 200
use FILL  FILL_13_1_0
timestamp 1556798218
transform -1 0 3224 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1556798218
transform -1 0 3240 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_2
timestamp 1556798218
transform -1 0 3256 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_296
timestamp 1556798218
transform -1 0 3448 0 1 2610
box 0 0 192 200
use AOI21X1  AOI21X1_72
timestamp 1556798218
transform -1 0 3512 0 1 2610
box 0 0 64 200
use INVX1  INVX1_499
timestamp 1556798218
transform -1 0 3544 0 1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_428
timestamp 1556798218
transform -1 0 3592 0 1 2610
box 0 0 48 200
use XNOR2X1  XNOR2X1_67
timestamp 1556798218
transform -1 0 3704 0 1 2610
box 0 0 112 200
use AOI22X1  AOI22X1_147
timestamp 1556798218
transform -1 0 3784 0 1 2610
box 0 0 80 200
use NAND2X1  NAND2X1_432
timestamp 1556798218
transform 1 0 3784 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_431
timestamp 1556798218
transform -1 0 3880 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_357
timestamp 1556798218
transform 1 0 3880 0 1 2610
box 0 0 192 200
use CLKBUF1  CLKBUF1_47
timestamp 1556798218
transform -1 0 4216 0 1 2610
box 0 0 144 200
use OAI21X1  OAI21X1_168
timestamp 1556798218
transform 1 0 4216 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_175
timestamp 1556798218
transform 1 0 4280 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_176
timestamp 1556798218
transform -1 0 4376 0 1 2610
box 0 0 48 200
use AOI22X1  AOI22X1_55
timestamp 1556798218
transform 1 0 4376 0 1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_71
timestamp 1556798218
transform 1 0 4456 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_14
timestamp 1556798218
transform 1 0 4504 0 1 2610
box 0 0 48 200
use INVX1  INVX1_176
timestamp 1556798218
transform 1 0 4552 0 1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_210
timestamp 1556798218
transform 1 0 4584 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_209
timestamp 1556798218
transform 1 0 4632 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_123
timestamp 1556798218
transform -1 0 4744 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_7
timestamp 1556798218
transform -1 0 4792 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_13
timestamp 1556798218
transform -1 0 4840 0 1 2610
box 0 0 48 200
use FILL  FILL_13_2_0
timestamp 1556798218
transform -1 0 4856 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1556798218
transform -1 0 4872 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_2
timestamp 1556798218
transform -1 0 4888 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_327
timestamp 1556798218
transform -1 0 5080 0 1 2610
box 0 0 192 200
use INVX1  INVX1_557
timestamp 1556798218
transform 1 0 5080 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_496
timestamp 1556798218
transform 1 0 5112 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_162
timestamp 1556798218
transform 1 0 5176 0 1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_218
timestamp 1556798218
transform 1 0 5256 0 1 2610
box 0 0 48 200
use AOI22X1  AOI22X1_163
timestamp 1556798218
transform -1 0 5384 0 1 2610
box 0 0 80 200
use NAND2X1  NAND2X1_478
timestamp 1556798218
transform 1 0 5384 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_477
timestamp 1556798218
transform 1 0 5432 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_474
timestamp 1556798218
transform -1 0 5528 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_127
timestamp 1556798218
transform -1 0 5592 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_491
timestamp 1556798218
transform 1 0 5592 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_492
timestamp 1556798218
transform -1 0 5720 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_6
timestamp 1556798218
transform 1 0 5720 0 1 2610
box 0 0 48 200
use INVX1  INVX1_256
timestamp 1556798218
transform 1 0 5768 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_236
timestamp 1556798218
transform 1 0 5800 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_77
timestamp 1556798218
transform 1 0 5864 0 1 2610
box 0 0 80 200
use AND2X2  AND2X2_65
timestamp 1556798218
transform -1 0 6008 0 1 2610
box 0 0 64 200
use INVX1  INVX1_255
timestamp 1556798218
transform 1 0 6008 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_234
timestamp 1556798218
transform 1 0 6040 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_233
timestamp 1556798218
transform -1 0 6168 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_154
timestamp 1556798218
transform -1 0 6360 0 1 2610
box 0 0 192 200
use FILL  FILL_13_3_0
timestamp 1556798218
transform 1 0 6360 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_1
timestamp 1556798218
transform 1 0 6376 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_2
timestamp 1556798218
transform 1 0 6392 0 1 2610
box 0 0 16 200
use XNOR2X1  XNOR2X1_32
timestamp 1556798218
transform 1 0 6408 0 1 2610
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_156
timestamp 1556798218
transform -1 0 6712 0 1 2610
box 0 0 192 200
use AND2X2  AND2X2_22
timestamp 1556798218
transform 1 0 6712 0 1 2610
box 0 0 64 200
use CLKBUF1  CLKBUF1_13
timestamp 1556798218
transform -1 0 6920 0 1 2610
box 0 0 144 200
use AND2X2  AND2X2_9
timestamp 1556798218
transform 1 0 6920 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_180
timestamp 1556798218
transform -1 0 7176 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_48
timestamp 1556798218
transform 1 0 7176 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_31
timestamp 1556798218
transform -1 0 7288 0 1 2610
box 0 0 64 200
use INVX1  INVX1_34
timestamp 1556798218
transform -1 0 7320 0 1 2610
box 0 0 32 200
use AOI22X1  AOI22X1_11
timestamp 1556798218
transform -1 0 7400 0 1 2610
box 0 0 80 200
use AOI22X1  AOI22X1_14
timestamp 1556798218
transform -1 0 7480 0 1 2610
box 0 0 80 200
use AOI22X1  AOI22X1_8
timestamp 1556798218
transform -1 0 7560 0 1 2610
box 0 0 80 200
use NAND2X1  NAND2X1_53
timestamp 1556798218
transform -1 0 7608 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1556798218
transform 1 0 7608 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_36
timestamp 1556798218
transform -1 0 7864 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_56
timestamp 1556798218
transform -1 0 7912 0 1 2610
box 0 0 48 200
use INVX1  INVX1_277
timestamp 1556798218
transform 1 0 7912 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_40
timestamp 1556798218
transform 1 0 7944 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_59
timestamp 1556798218
transform -1 0 8056 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_263
timestamp 1556798218
transform -1 0 8104 0 1 2610
box 0 0 48 200
use INVX1  INVX1_196
timestamp 1556798218
transform -1 0 8136 0 1 2610
box 0 0 32 200
use FILL  FILL_14_1
timestamp 1556798218
transform 1 0 8136 0 1 2610
box 0 0 16 200
use FILL  FILL_14_2
timestamp 1556798218
transform 1 0 8152 0 1 2610
box 0 0 16 200
use CLKBUF1  CLKBUF1_50
timestamp 1556798218
transform -1 0 152 0 -1 2610
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_365
timestamp 1556798218
transform -1 0 344 0 -1 2610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_232
timestamp 1556798218
transform -1 0 536 0 -1 2610
box 0 0 192 200
use INVX1  INVX1_619
timestamp 1556798218
transform 1 0 536 0 -1 2610
box 0 0 32 200
use BUFX2  BUFX2_8
timestamp 1556798218
transform -1 0 616 0 -1 2610
box 0 0 48 200
use CLKBUF1  CLKBUF1_39
timestamp 1556798218
transform 1 0 616 0 -1 2610
box 0 0 144 200
use INVX1  INVX1_385
timestamp 1556798218
transform -1 0 792 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_351
timestamp 1556798218
transform 1 0 792 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_343
timestamp 1556798218
transform -1 0 904 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_384
timestamp 1556798218
transform -1 0 936 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_347
timestamp 1556798218
transform -1 0 1000 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_386
timestamp 1556798218
transform 1 0 1000 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_348
timestamp 1556798218
transform -1 0 1096 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_114
timestamp 1556798218
transform -1 0 1176 0 -1 2610
box 0 0 80 200
use BUFX2  BUFX2_37
timestamp 1556798218
transform 1 0 1176 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_379
timestamp 1556798218
transform 1 0 1224 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_340
timestamp 1556798218
transform -1 0 1304 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_341
timestamp 1556798218
transform -1 0 1352 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_144
timestamp 1556798218
transform -1 0 1400 0 -1 2610
box 0 0 48 200
use AOI22X1  AOI22X1_113
timestamp 1556798218
transform -1 0 1480 0 -1 2610
box 0 0 80 200
use INVX1  INVX1_380
timestamp 1556798218
transform 1 0 1480 0 -1 2610
box 0 0 32 200
use INVX1  INVX1_378
timestamp 1556798218
transform 1 0 1512 0 -1 2610
box 0 0 32 200
use AOI22X1  AOI22X1_112
timestamp 1556798218
transform -1 0 1624 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_342
timestamp 1556798218
transform -1 0 1688 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_341
timestamp 1556798218
transform -1 0 1752 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_0_0
timestamp 1556798218
transform -1 0 1768 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1556798218
transform -1 0 1784 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_2
timestamp 1556798218
transform -1 0 1800 0 -1 2610
box 0 0 16 200
use NAND3X1  NAND3X1_116
timestamp 1556798218
transform -1 0 1864 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_117
timestamp 1556798218
transform -1 0 1928 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_345
timestamp 1556798218
transform 1 0 1928 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_143
timestamp 1556798218
transform 1 0 1992 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_376
timestamp 1556798218
transform -1 0 2072 0 -1 2610
box 0 0 32 200
use CLKBUF1  CLKBUF1_1
timestamp 1556798218
transform 1 0 2072 0 -1 2610
box 0 0 144 200
use NOR2X1  NOR2X1_123
timestamp 1556798218
transform 1 0 2216 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_124
timestamp 1556798218
transform 1 0 2264 0 -1 2610
box 0 0 48 200
use AND2X2  AND2X2_80
timestamp 1556798218
transform -1 0 2376 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1556798218
transform -1 0 2440 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_102
timestamp 1556798218
transform -1 0 2472 0 -1 2610
box 0 0 32 200
use AND2X2  AND2X2_78
timestamp 1556798218
transform 1 0 2472 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_119
timestamp 1556798218
transform -1 0 2584 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_96
timestamp 1556798218
transform 1 0 2584 0 -1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_46
timestamp 1556798218
transform -1 0 2664 0 -1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_68
timestamp 1556798218
transform -1 0 2856 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_429
timestamp 1556798218
transform 1 0 2856 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_447
timestamp 1556798218
transform 1 0 2904 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_444
timestamp 1556798218
transform 1 0 2968 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_443
timestamp 1556798218
transform -1 0 3096 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_498
timestamp 1556798218
transform 1 0 3096 0 -1 2610
box 0 0 32 200
use INVX1  INVX1_497
timestamp 1556798218
transform -1 0 3160 0 -1 2610
box 0 0 32 200
use AOI22X1  AOI22X1_146
timestamp 1556798218
transform 1 0 3160 0 -1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_150
timestamp 1556798218
transform 1 0 3240 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_1_0
timestamp 1556798218
transform -1 0 3320 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1556798218
transform -1 0 3336 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_2
timestamp 1556798218
transform -1 0 3352 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_430
timestamp 1556798218
transform -1 0 3400 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_496
timestamp 1556798218
transform -1 0 3432 0 -1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_190
timestamp 1556798218
transform -1 0 3480 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_445
timestamp 1556798218
transform 1 0 3480 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_446
timestamp 1556798218
transform -1 0 3608 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_294
timestamp 1556798218
transform 1 0 3608 0 -1 2610
box 0 0 192 200
use INVX1  INVX1_500
timestamp 1556798218
transform -1 0 3832 0 -1 2610
box 0 0 32 200
use AND2X2  AND2X2_113
timestamp 1556798218
transform -1 0 3896 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_111
timestamp 1556798218
transform -1 0 4088 0 -1 2610
box 0 0 192 200
use AND2X2  AND2X2_128
timestamp 1556798218
transform 1 0 4088 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_179
timestamp 1556798218
transform 1 0 4152 0 -1 2610
box 0 0 32 200
use AOI22X1  AOI22X1_165
timestamp 1556798218
transform 1 0 4184 0 -1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_220
timestamp 1556798218
transform -1 0 4312 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_482
timestamp 1556798218
transform 1 0 4312 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_483
timestamp 1556798218
transform -1 0 4408 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_561
timestamp 1556798218
transform -1 0 4440 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_479
timestamp 1556798218
transform 1 0 4440 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_168
timestamp 1556798218
transform -1 0 4552 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_563
timestamp 1556798218
transform 1 0 4552 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_467
timestamp 1556798218
transform 1 0 4584 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_500
timestamp 1556798218
transform 1 0 4632 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_330
timestamp 1556798218
transform 1 0 4696 0 -1 2610
box 0 0 192 200
use FILL  FILL_12_2_0
timestamp 1556798218
transform 1 0 4888 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1556798218
transform 1 0 4904 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_2
timestamp 1556798218
transform 1 0 4920 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_326
timestamp 1556798218
transform 1 0 4936 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_475
timestamp 1556798218
transform 1 0 5128 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_552
timestamp 1556798218
transform -1 0 5208 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_476
timestamp 1556798218
transform 1 0 5208 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_493
timestamp 1556798218
transform 1 0 5256 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_494
timestamp 1556798218
transform -1 0 5384 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_556
timestamp 1556798218
transform -1 0 5416 0 -1 2610
box 0 0 32 200
use BUFX2  BUFX2_97
timestamp 1556798218
transform -1 0 5464 0 -1 2610
box 0 0 48 200
use BUFX2  BUFX2_95
timestamp 1556798218
transform 1 0 5464 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_11
timestamp 1556798218
transform 1 0 5512 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_239
timestamp 1556798218
transform 1 0 5560 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_238
timestamp 1556798218
transform -1 0 5656 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_253
timestamp 1556798218
transform 1 0 5656 0 -1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_95
timestamp 1556798218
transform -1 0 5736 0 -1 2610
box 0 0 48 200
use AOI22X1  AOI22X1_76
timestamp 1556798218
transform -1 0 5816 0 -1 2610
box 0 0 80 200
use INVX1  INVX1_251
timestamp 1556798218
transform -1 0 5848 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_237
timestamp 1556798218
transform 1 0 5848 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_80
timestamp 1556798218
transform -1 0 5960 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_231
timestamp 1556798218
transform 1 0 5960 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_235
timestamp 1556798218
transform 1 0 6024 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_232
timestamp 1556798218
transform -1 0 6136 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_252
timestamp 1556798218
transform 1 0 6136 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_236
timestamp 1556798218
transform -1 0 6216 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_254
timestamp 1556798218
transform -1 0 6248 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_235
timestamp 1556798218
transform 1 0 6248 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_37
timestamp 1556798218
transform -1 0 6376 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_3_0
timestamp 1556798218
transform -1 0 6392 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_1
timestamp 1556798218
transform -1 0 6408 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_2
timestamp 1556798218
transform -1 0 6424 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_157
timestamp 1556798218
transform -1 0 6616 0 -1 2610
box 0 0 192 200
use BUFX2  BUFX2_69
timestamp 1556798218
transform 1 0 6616 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_412
timestamp 1556798218
transform -1 0 6728 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_459
timestamp 1556798218
transform -1 0 6760 0 -1 2610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_271
timestamp 1556798218
transform 1 0 6760 0 -1 2610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1556798218
transform -1 0 7144 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_51
timestamp 1556798218
transform 1 0 7144 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_34
timestamp 1556798218
transform -1 0 7256 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_37
timestamp 1556798218
transform -1 0 7288 0 -1 2610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1556798218
transform 1 0 7288 0 -1 2610
box 0 0 192 200
use NAND3X1  NAND3X1_16
timestamp 1556798218
transform 1 0 7480 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_4
timestamp 1556798218
transform 1 0 7544 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_28
timestamp 1556798218
transform 1 0 7608 0 -1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_22
timestamp 1556798218
transform 1 0 7640 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_35
timestamp 1556798218
transform 1 0 7688 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_52
timestamp 1556798218
transform -1 0 7800 0 -1 2610
box 0 0 48 200
use AND2X2  AND2X2_24
timestamp 1556798218
transform 1 0 7800 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1556798218
transform 1 0 7864 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1556798218
transform 1 0 7928 0 -1 2610
box 0 0 192 200
use FILL  FILL_13_1
timestamp 1556798218
transform -1 0 8136 0 -1 2610
box 0 0 16 200
use FILL  FILL_13_2
timestamp 1556798218
transform -1 0 8152 0 -1 2610
box 0 0 16 200
use FILL  FILL_13_3
timestamp 1556798218
transform -1 0 8168 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_364
timestamp 1556798218
transform 1 0 8 0 1 2210
box 0 0 192 200
use INVX1  INVX1_618
timestamp 1556798218
transform -1 0 232 0 1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_523
timestamp 1556798218
transform 1 0 232 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_185
timestamp 1556798218
transform 1 0 280 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_184
timestamp 1556798218
transform 1 0 344 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_524
timestamp 1556798218
transform 1 0 408 0 1 2210
box 0 0 48 200
use INVX1  INVX1_615
timestamp 1556798218
transform -1 0 488 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_547
timestamp 1556798218
transform 1 0 488 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_548
timestamp 1556798218
transform 1 0 552 0 1 2210
box 0 0 64 200
use INVX1  INVX1_617
timestamp 1556798218
transform -1 0 648 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_362
timestamp 1556798218
transform -1 0 840 0 1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_233
timestamp 1556798218
transform -1 0 1032 0 1 2210
box 0 0 192 200
use NAND3X1  NAND3X1_119
timestamp 1556798218
transform 1 0 1032 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_118
timestamp 1556798218
transform -1 0 1160 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_349
timestamp 1556798218
transform 1 0 1160 0 1 2210
box 0 0 64 200
use INVX1  INVX1_387
timestamp 1556798218
transform -1 0 1256 0 1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_342
timestamp 1556798218
transform -1 0 1304 0 1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_146
timestamp 1556798218
transform -1 0 1352 0 1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_115
timestamp 1556798218
transform -1 0 1432 0 1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_346
timestamp 1556798218
transform -1 0 1480 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_334
timestamp 1556798218
transform 1 0 1480 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_352
timestamp 1556798218
transform -1 0 1592 0 1 2210
box 0 0 64 200
use INVX1  INVX1_389
timestamp 1556798218
transform -1 0 1624 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_231
timestamp 1556798218
transform 1 0 1624 0 1 2210
box 0 0 192 200
use FILL  FILL_11_0_0
timestamp 1556798218
transform -1 0 1832 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1556798218
transform -1 0 1848 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_2
timestamp 1556798218
transform -1 0 1864 0 1 2210
box 0 0 16 200
use NOR2X1  NOR2X1_122
timestamp 1556798218
transform -1 0 1912 0 1 2210
box 0 0 48 200
use AND2X2  AND2X2_79
timestamp 1556798218
transform -1 0 1976 0 1 2210
box 0 0 64 200
use INVX1  INVX1_382
timestamp 1556798218
transform 1 0 1976 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_346
timestamp 1556798218
transform 1 0 2008 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_121
timestamp 1556798218
transform -1 0 2120 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_229
timestamp 1556798218
transform -1 0 2312 0 1 2210
box 0 0 192 200
use NOR2X1  NOR2X1_52
timestamp 1556798218
transform 1 0 2312 0 1 2210
box 0 0 48 200
use INVX1  INVX1_117
timestamp 1556798218
transform -1 0 2392 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_69
timestamp 1556798218
transform 1 0 2392 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_109
timestamp 1556798218
transform 1 0 2584 0 1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_32
timestamp 1556798218
transform 1 0 2632 0 1 2210
box 0 0 80 200
use INVX1  INVX1_98
timestamp 1556798218
transform 1 0 2712 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_95
timestamp 1556798218
transform 1 0 2744 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_96
timestamp 1556798218
transform -1 0 2872 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_37
timestamp 1556798218
transform -1 0 2936 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_99
timestamp 1556798218
transform -1 0 3000 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_110
timestamp 1556798218
transform -1 0 3048 0 1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_15
timestamp 1556798218
transform -1 0 3112 0 1 2210
box 0 0 64 200
use BUFX2  BUFX2_71
timestamp 1556798218
transform -1 0 3160 0 1 2210
box 0 0 48 200
use INVX1  INVX1_495
timestamp 1556798218
transform 1 0 3160 0 1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_189
timestamp 1556798218
transform -1 0 3240 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_151
timestamp 1556798218
transform 1 0 3240 0 1 2210
box 0 0 64 200
use FILL  FILL_11_1_0
timestamp 1556798218
transform 1 0 3304 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1556798218
transform 1 0 3320 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_2
timestamp 1556798218
transform 1 0 3336 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_297
timestamp 1556798218
transform 1 0 3352 0 1 2210
box 0 0 192 200
use CLKBUF1  CLKBUF1_23
timestamp 1556798218
transform -1 0 3688 0 1 2210
box 0 0 144 200
use BUFX2  BUFX2_130
timestamp 1556798218
transform -1 0 3736 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_334
timestamp 1556798218
transform 1 0 3736 0 1 2210
box 0 0 192 200
use BUFX2  BUFX2_132
timestamp 1556798218
transform -1 0 3976 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_506
timestamp 1556798218
transform -1 0 4040 0 1 2210
box 0 0 64 200
use INVX1  INVX1_570
timestamp 1556798218
transform -1 0 4072 0 1 2210
box 0 0 32 200
use AND2X2  AND2X2_129
timestamp 1556798218
transform 1 0 4072 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_333
timestamp 1556798218
transform -1 0 4328 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_502
timestamp 1556798218
transform -1 0 4392 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_164
timestamp 1556798218
transform -1 0 4472 0 1 2210
box 0 0 80 200
use INVX1  INVX1_562
timestamp 1556798218
transform 1 0 4472 0 1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_481
timestamp 1556798218
transform -1 0 4552 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_169
timestamp 1556798218
transform 1 0 4552 0 1 2210
box 0 0 64 200
use INVX1  INVX1_560
timestamp 1556798218
transform 1 0 4616 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_497
timestamp 1556798218
transform 1 0 4648 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_498
timestamp 1556798218
transform -1 0 4776 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_499
timestamp 1556798218
transform -1 0 4840 0 1 2210
box 0 0 64 200
use FILL  FILL_11_2_0
timestamp 1556798218
transform -1 0 4856 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1556798218
transform -1 0 4872 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_2
timestamp 1556798218
transform -1 0 4888 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_501
timestamp 1556798218
transform -1 0 4952 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_81
timestamp 1556798218
transform -1 0 5016 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_480
timestamp 1556798218
transform -1 0 5064 0 1 2210
box 0 0 48 200
use INVX1  INVX1_559
timestamp 1556798218
transform -1 0 5096 0 1 2210
box 0 0 32 200
use XNOR2X1  XNOR2X1_76
timestamp 1556798218
transform -1 0 5208 0 1 2210
box 0 0 112 200
use BUFX2  BUFX2_125
timestamp 1556798218
transform -1 0 5256 0 1 2210
box 0 0 48 200
use CLKBUF1  CLKBUF1_17
timestamp 1556798218
transform 1 0 5256 0 1 2210
box 0 0 144 200
use NAND2X1  NAND2X1_380
timestamp 1556798218
transform 1 0 5400 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_392
timestamp 1556798218
transform 1 0 5448 0 1 2210
box 0 0 64 200
use INVX1  INVX1_437
timestamp 1556798218
transform -1 0 5544 0 1 2210
box 0 0 32 200
use AND2X2  AND2X2_101
timestamp 1556798218
transform -1 0 5608 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_391
timestamp 1556798218
transform -1 0 5672 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_128
timestamp 1556798218
transform -1 0 5752 0 1 2210
box 0 0 80 200
use BUFX2  BUFX2_96
timestamp 1556798218
transform 1 0 5752 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_132
timestamp 1556798218
transform -1 0 5864 0 1 2210
box 0 0 64 200
use INVX1  INVX1_435
timestamp 1556798218
transform -1 0 5896 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_389
timestamp 1556798218
transform 1 0 5896 0 1 2210
box 0 0 64 200
use INVX1  INVX1_434
timestamp 1556798218
transform 1 0 5960 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_393
timestamp 1556798218
transform 1 0 5992 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_133
timestamp 1556798218
transform 1 0 6056 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_390
timestamp 1556798218
transform -1 0 6184 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_165
timestamp 1556798218
transform 1 0 6184 0 1 2210
box 0 0 48 200
use INVX1  INVX1_432
timestamp 1556798218
transform -1 0 6264 0 1 2210
box 0 0 32 200
use NAND3X1  NAND3X1_81
timestamp 1556798218
transform -1 0 6328 0 1 2210
box 0 0 64 200
use INVX1  INVX1_250
timestamp 1556798218
transform 1 0 6328 0 1 2210
box 0 0 32 200
use FILL  FILL_11_3_0
timestamp 1556798218
transform -1 0 6376 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_1
timestamp 1556798218
transform -1 0 6392 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_2
timestamp 1556798218
transform -1 0 6408 0 1 2210
box 0 0 16 200
use NOR2X1  NOR2X1_94
timestamp 1556798218
transform -1 0 6456 0 1 2210
box 0 0 48 200
use INVX1  INVX1_456
timestamp 1556798218
transform 1 0 6456 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_272
timestamp 1556798218
transform 1 0 6488 0 1 2210
box 0 0 192 200
use AOI22X1  AOI22X1_134
timestamp 1556798218
transform -1 0 6760 0 1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_399
timestamp 1556798218
transform 1 0 6760 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_396
timestamp 1556798218
transform -1 0 6856 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_398
timestamp 1556798218
transform -1 0 6904 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_49
timestamp 1556798218
transform 1 0 6904 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_32
timestamp 1556798218
transform -1 0 7016 0 1 2210
box 0 0 64 200
use INVX1  INVX1_35
timestamp 1556798218
transform -1 0 7048 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1556798218
transform 1 0 7048 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_46
timestamp 1556798218
transform -1 0 7288 0 1 2210
box 0 0 48 200
use INVX1  INVX1_26
timestamp 1556798218
transform 1 0 7288 0 1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_20
timestamp 1556798218
transform -1 0 7368 0 1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_23
timestamp 1556798218
transform 1 0 7368 0 1 2210
box 0 0 48 200
use INVX1  INVX1_27
timestamp 1556798218
transform 1 0 7416 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_37
timestamp 1556798218
transform 1 0 7448 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_21
timestamp 1556798218
transform 1 0 7512 0 1 2210
box 0 0 48 200
use INVX1  INVX1_29
timestamp 1556798218
transform -1 0 7592 0 1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_44
timestamp 1556798218
transform -1 0 7640 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_26
timestamp 1556798218
transform 1 0 7640 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_27
timestamp 1556798218
transform -1 0 7768 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_15
timestamp 1556798218
transform 1 0 7768 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1556798218
transform 1 0 7832 0 1 2210
box 0 0 64 200
use INVX1  INVX1_31
timestamp 1556798218
transform -1 0 7928 0 1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1556798218
transform 1 0 7928 0 1 2210
box 0 0 192 200
use FILL  FILL_12_1
timestamp 1556798218
transform 1 0 8120 0 1 2210
box 0 0 16 200
use FILL  FILL_12_2
timestamp 1556798218
transform 1 0 8136 0 1 2210
box 0 0 16 200
use FILL  FILL_12_3
timestamp 1556798218
transform 1 0 8152 0 1 2210
box 0 0 16 200
use XNOR2X1  XNOR2X1_84
timestamp 1556798218
transform 1 0 8 0 -1 2210
box 0 0 112 200
use AOI21X1  AOI21X1_89
timestamp 1556798218
transform 1 0 120 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_616
timestamp 1556798218
transform 1 0 184 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_549
timestamp 1556798218
transform 1 0 216 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_546
timestamp 1556798218
transform 1 0 280 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_545
timestamp 1556798218
transform -1 0 408 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_180
timestamp 1556798218
transform -1 0 488 0 -1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_522
timestamp 1556798218
transform 1 0 488 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_526
timestamp 1556798218
transform 1 0 536 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_181
timestamp 1556798218
transform 1 0 584 0 -1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_525
timestamp 1556798218
transform -1 0 712 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_242
timestamp 1556798218
transform 1 0 712 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_241
timestamp 1556798218
transform 1 0 760 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_230
timestamp 1556798218
transform 1 0 952 0 -1 2210
box 0 0 192 200
use BUFX2  BUFX2_79
timestamp 1556798218
transform 1 0 1144 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_350
timestamp 1556798218
transform -1 0 1256 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_388
timestamp 1556798218
transform -1 0 1288 0 -1 2210
box 0 0 32 200
use AND2X2  AND2X2_91
timestamp 1556798218
transform 1 0 1288 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_345
timestamp 1556798218
transform 1 0 1352 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_335
timestamp 1556798218
transform 1 0 1400 0 -1 2210
box 0 0 48 200
use NOR3X1  NOR3X1_3
timestamp 1556798218
transform 1 0 1448 0 -1 2210
box 0 0 128 200
use NOR2X1  NOR2X1_138
timestamp 1556798218
transform 1 0 1576 0 -1 2210
box 0 0 48 200
use AND2X2  AND2X2_87
timestamp 1556798218
transform -1 0 1688 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_137
timestamp 1556798218
transform 1 0 1688 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_0_0
timestamp 1556798218
transform 1 0 1736 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1556798218
transform 1 0 1752 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_2
timestamp 1556798218
transform 1 0 1768 0 -1 2210
box 0 0 16 200
use AND2X2  AND2X2_89
timestamp 1556798218
transform 1 0 1784 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_141
timestamp 1556798218
transform 1 0 1848 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_142
timestamp 1556798218
transform 1 0 1896 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_227
timestamp 1556798218
transform -1 0 2136 0 -1 2210
box 0 0 192 200
use NOR3X1  NOR3X1_2
timestamp 1556798218
transform 1 0 2136 0 -1 2210
box 0 0 128 200
use BUFX2  BUFX2_80
timestamp 1556798218
transform 1 0 2264 0 -1 2210
box 0 0 48 200
use BUFX2  BUFX2_104
timestamp 1556798218
transform 1 0 2312 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_66
timestamp 1556798218
transform 1 0 2360 0 -1 2210
box 0 0 192 200
use AOI22X1  AOI22X1_33
timestamp 1556798218
transform -1 0 2632 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_98
timestamp 1556798218
transform 1 0 2632 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_47
timestamp 1556798218
transform 1 0 2696 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_97
timestamp 1556798218
transform -1 0 2808 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_113
timestamp 1556798218
transform -1 0 2856 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_111
timestamp 1556798218
transform -1 0 2904 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_36
timestamp 1556798218
transform 1 0 2904 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_99
timestamp 1556798218
transform -1 0 3000 0 -1 2210
box 0 0 32 200
use INVX1  INVX1_97
timestamp 1556798218
transform -1 0 3032 0 -1 2210
box 0 0 32 200
use XNOR2X1  XNOR2X1_10
timestamp 1556798218
transform -1 0 3144 0 -1 2210
box 0 0 112 200
use INVX1  INVX1_100
timestamp 1556798218
transform -1 0 3176 0 -1 2210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_253
timestamp 1556798218
transform -1 0 3368 0 -1 2210
box 0 0 192 200
use FILL  FILL_10_1_0
timestamp 1556798218
transform 1 0 3368 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1556798218
transform 1 0 3384 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_2
timestamp 1556798218
transform 1 0 3400 0 -1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_129
timestamp 1556798218
transform 1 0 3416 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_302
timestamp 1556798218
transform -1 0 3528 0 -1 2210
box 0 0 48 200
use XNOR2X1  XNOR2X1_77
timestamp 1556798218
transform 1 0 3528 0 -1 2210
box 0 0 112 200
use AOI21X1  AOI21X1_82
timestamp 1556798218
transform 1 0 3640 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_565
timestamp 1556798218
transform 1 0 3704 0 -1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_221
timestamp 1556798218
transform -1 0 3784 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_507
timestamp 1556798218
transform -1 0 3848 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_485
timestamp 1556798218
transform 1 0 3848 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_566
timestamp 1556798218
transform 1 0 3896 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_505
timestamp 1556798218
transform 1 0 3928 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_484
timestamp 1556798218
transform -1 0 4040 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_567
timestamp 1556798218
transform -1 0 4072 0 -1 2210
box 0 0 32 200
use BUFX2  BUFX2_123
timestamp 1556798218
transform -1 0 4120 0 -1 2210
box 0 0 48 200
use CLKBUF1  CLKBUF1_42
timestamp 1556798218
transform 1 0 4120 0 -1 2210
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_331
timestamp 1556798218
transform 1 0 4264 0 -1 2210
box 0 0 192 200
use INVX1  INVX1_564
timestamp 1556798218
transform -1 0 4488 0 -1 2210
box 0 0 32 200
use BUFX2  BUFX2_98
timestamp 1556798218
transform 1 0 4488 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_219
timestamp 1556798218
transform 1 0 4536 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_332
timestamp 1556798218
transform -1 0 4776 0 -1 2210
box 0 0 192 200
use FILL  FILL_10_2_0
timestamp 1556798218
transform -1 0 4792 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1556798218
transform -1 0 4808 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_2
timestamp 1556798218
transform -1 0 4824 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_285
timestamp 1556798218
transform -1 0 5016 0 -1 2210
box 0 0 192 200
use NAND3X1  NAND3X1_145
timestamp 1556798218
transform 1 0 5016 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_476
timestamp 1556798218
transform -1 0 5112 0 -1 2210
box 0 0 32 200
use BUFX2  BUFX2_101
timestamp 1556798218
transform 1 0 5112 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_258
timestamp 1556798218
transform 1 0 5160 0 -1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_383
timestamp 1556798218
transform -1 0 5400 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_384
timestamp 1556798218
transform -1 0 5448 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_129
timestamp 1556798218
transform 1 0 5448 0 -1 2210
box 0 0 80 200
use NOR2X1  NOR2X1_166
timestamp 1556798218
transform 1 0 5528 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_436
timestamp 1556798218
transform 1 0 5576 0 -1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_382
timestamp 1556798218
transform -1 0 5656 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_433
timestamp 1556798218
transform -1 0 5688 0 -1 2210
box 0 0 32 200
use XNOR2X1  XNOR2X1_58
timestamp 1556798218
transform -1 0 5800 0 -1 2210
box 0 0 112 200
use AOI21X1  AOI21X1_63
timestamp 1556798218
transform 1 0 5800 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_381
timestamp 1556798218
transform 1 0 5864 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_261
timestamp 1556798218
transform -1 0 6104 0 -1 2210
box 0 0 192 200
use XNOR2X1  XNOR2X1_61
timestamp 1556798218
transform -1 0 6216 0 -1 2210
box 0 0 112 200
use AND2X2  AND2X2_63
timestamp 1556798218
transform 1 0 6216 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_248
timestamp 1556798218
transform 1 0 6280 0 -1 2210
box 0 0 32 200
use AOI21X1  AOI21X1_66
timestamp 1556798218
transform 1 0 6312 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_3_0
timestamp 1556798218
transform -1 0 6392 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_1
timestamp 1556798218
transform -1 0 6408 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_2
timestamp 1556798218
transform -1 0 6424 0 -1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_138
timestamp 1556798218
transform -1 0 6488 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_397
timestamp 1556798218
transform 1 0 6488 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_172
timestamp 1556798218
transform -1 0 6584 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_135
timestamp 1556798218
transform -1 0 6664 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_407
timestamp 1556798218
transform 1 0 6664 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_408
timestamp 1556798218
transform -1 0 6792 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_411
timestamp 1556798218
transform 1 0 6792 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_139
timestamp 1556798218
transform -1 0 6920 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_453
timestamp 1556798218
transform 1 0 6920 0 -1 2210
box 0 0 32 200
use NOR2X1  NOR2X1_171
timestamp 1556798218
transform -1 0 7000 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_50
timestamp 1556798218
transform 1 0 7000 0 -1 2210
box 0 0 48 200
use AOI22X1  AOI22X1_12
timestamp 1556798218
transform -1 0 7128 0 -1 2210
box 0 0 80 200
use AOI22X1  AOI22X1_13
timestamp 1556798218
transform -1 0 7208 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_29
timestamp 1556798218
transform 1 0 7208 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_32
timestamp 1556798218
transform -1 0 7304 0 -1 2210
box 0 0 32 200
use AOI22X1  AOI22X1_9
timestamp 1556798218
transform -1 0 7384 0 -1 2210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1556798218
transform -1 0 7576 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1556798218
transform -1 0 7768 0 -1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_58
timestamp 1556798218
transform -1 0 7816 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_42
timestamp 1556798218
transform 1 0 7816 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1556798218
transform 1 0 7880 0 -1 2210
box 0 0 192 200
use BUFX2  BUFX2_142
timestamp 1556798218
transform 1 0 8072 0 -1 2210
box 0 0 48 200
use FILL  FILL_11_1
timestamp 1556798218
transform -1 0 8136 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1556798218
transform -1 0 8152 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_3
timestamp 1556798218
transform -1 0 8168 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_105
timestamp 1556798218
transform 1 0 8 0 1 1810
box 0 0 192 200
use AND2X2  AND2X2_20
timestamp 1556798218
transform 1 0 200 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_241
timestamp 1556798218
transform 1 0 264 0 1 1810
box 0 0 48 200
use INVX1  INVX1_614
timestamp 1556798218
transform -1 0 344 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_550
timestamp 1556798218
transform -1 0 408 0 1 1810
box 0 0 64 200
use INVX1  INVX1_620
timestamp 1556798218
transform -1 0 440 0 1 1810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_363
timestamp 1556798218
transform 1 0 440 0 1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_123
timestamp 1556798218
transform 1 0 632 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_360
timestamp 1556798218
transform 1 0 696 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_359
timestamp 1556798218
transform -1 0 824 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_122
timestamp 1556798218
transform 1 0 824 0 1 1810
box 0 0 64 200
use INVX1  INVX1_399
timestamp 1556798218
transform -1 0 920 0 1 1810
box 0 0 32 200
use INVX1  INVX1_400
timestamp 1556798218
transform -1 0 952 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_354
timestamp 1556798218
transform 1 0 952 0 1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_118
timestamp 1556798218
transform -1 0 1080 0 1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_150
timestamp 1556798218
transform -1 0 1128 0 1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_119
timestamp 1556798218
transform -1 0 1208 0 1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_364
timestamp 1556798218
transform -1 0 1272 0 1 1810
box 0 0 64 200
use INVX1  INVX1_403
timestamp 1556798218
transform -1 0 1304 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_85
timestamp 1556798218
transform -1 0 1368 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_93
timestamp 1556798218
transform -1 0 1432 0 1 1810
box 0 0 64 200
use BUFX2  BUFX2_120
timestamp 1556798218
transform -1 0 1480 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_239
timestamp 1556798218
transform -1 0 1672 0 1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_139
timestamp 1556798218
transform 1 0 1672 0 1 1810
box 0 0 48 200
use FILL  FILL_9_0_0
timestamp 1556798218
transform 1 0 1720 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1556798218
transform 1 0 1736 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_2
timestamp 1556798218
transform 1 0 1752 0 1 1810
box 0 0 16 200
use AND2X2  AND2X2_88
timestamp 1556798218
transform 1 0 1768 0 1 1810
box 0 0 64 200
use BUFX2  BUFX2_38
timestamp 1556798218
transform -1 0 1880 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_81
timestamp 1556798218
transform 1 0 1880 0 1 1810
box 0 0 192 200
use BUFX2  BUFX2_35
timestamp 1556798218
transform -1 0 2120 0 1 1810
box 0 0 48 200
use INVX1  INVX1_119
timestamp 1556798218
transform 1 0 2120 0 1 1810
box 0 0 32 200
use BUFX2  BUFX2_105
timestamp 1556798218
transform 1 0 2152 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_43
timestamp 1556798218
transform -1 0 2264 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1556798218
transform -1 0 2328 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_127
timestamp 1556798218
transform 1 0 2328 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_115
timestamp 1556798218
transform 1 0 2376 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_114
timestamp 1556798218
transform -1 0 2504 0 1 1810
box 0 0 64 200
use INVX1  INVX1_120
timestamp 1556798218
transform -1 0 2536 0 1 1810
box 0 0 32 200
use INVX1  INVX1_118
timestamp 1556798218
transform -1 0 2568 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_39
timestamp 1556798218
transform 1 0 2568 0 1 1810
box 0 0 64 200
use INVX1  INVX1_101
timestamp 1556798218
transform -1 0 2664 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_129
timestamp 1556798218
transform -1 0 2712 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_130
timestamp 1556798218
transform -1 0 2760 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_126
timestamp 1556798218
transform -1 0 2808 0 1 1810
box 0 0 48 200
use AND2X2  AND2X2_99
timestamp 1556798218
transform 1 0 2808 0 1 1810
box 0 0 64 200
use INVX1  INVX1_423
timestamp 1556798218
transform 1 0 2872 0 1 1810
box 0 0 32 200
use XNOR2X1  XNOR2X1_56
timestamp 1556798218
transform -1 0 3016 0 1 1810
box 0 0 112 200
use AOI21X1  AOI21X1_61
timestamp 1556798218
transform 1 0 3016 0 1 1810
box 0 0 64 200
use INVX1  INVX1_420
timestamp 1556798218
transform 1 0 3080 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_381
timestamp 1556798218
transform 1 0 3112 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_371
timestamp 1556798218
transform 1 0 3176 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_377
timestamp 1556798218
transform -1 0 3288 0 1 1810
box 0 0 64 200
use FILL  FILL_9_1_0
timestamp 1556798218
transform -1 0 3304 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1556798218
transform -1 0 3320 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_2
timestamp 1556798218
transform -1 0 3336 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_378
timestamp 1556798218
transform -1 0 3400 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_128
timestamp 1556798218
transform -1 0 3464 0 1 1810
box 0 0 64 200
use INVX1  INVX1_418
timestamp 1556798218
transform 1 0 3464 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_161
timestamp 1556798218
transform -1 0 3544 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_336
timestamp 1556798218
transform 1 0 3544 0 1 1810
box 0 0 192 200
use INVX1  INVX1_569
timestamp 1556798218
transform 1 0 3736 0 1 1810
box 0 0 32 200
use INVX1  INVX1_568
timestamp 1556798218
transform 1 0 3768 0 1 1810
box 0 0 32 200
use NAND3X1  NAND3X1_170
timestamp 1556798218
transform -1 0 3864 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_171
timestamp 1556798218
transform 1 0 3864 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_504
timestamp 1556798218
transform 1 0 3928 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_503
timestamp 1556798218
transform -1 0 4056 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_486
timestamp 1556798218
transform 1 0 4056 0 1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_166
timestamp 1556798218
transform -1 0 4184 0 1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_222
timestamp 1556798218
transform -1 0 4232 0 1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_167
timestamp 1556798218
transform -1 0 4312 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_488
timestamp 1556798218
transform 1 0 4312 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_487
timestamp 1556798218
transform -1 0 4408 0 1 1810
box 0 0 48 200
use AND2X2  AND2X2_50
timestamp 1556798218
transform -1 0 4472 0 1 1810
box 0 0 64 200
use INVX1  INVX1_466
timestamp 1556798218
transform -1 0 4504 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_178
timestamp 1556798218
transform -1 0 4552 0 1 1810
box 0 0 48 200
use INVX1  INVX1_558
timestamp 1556798218
transform 1 0 4552 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_107
timestamp 1556798218
transform -1 0 4648 0 1 1810
box 0 0 64 200
use XNOR2X1  XNOR2X1_64
timestamp 1556798218
transform -1 0 4760 0 1 1810
box 0 0 112 200
use INVX1  INVX1_474
timestamp 1556798218
transform 1 0 4760 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_183
timestamp 1556798218
transform -1 0 4840 0 1 1810
box 0 0 48 200
use FILL  FILL_9_2_0
timestamp 1556798218
transform 1 0 4840 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1556798218
transform 1 0 4856 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_2
timestamp 1556798218
transform 1 0 4872 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_69
timestamp 1556798218
transform 1 0 4888 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_429
timestamp 1556798218
transform -1 0 5016 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_144
timestamp 1556798218
transform -1 0 5080 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_425
timestamp 1556798218
transform -1 0 5144 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_426
timestamp 1556798218
transform -1 0 5208 0 1 1810
box 0 0 64 200
use INVX1  INVX1_475
timestamp 1556798218
transform -1 0 5240 0 1 1810
box 0 0 32 200
use INVX1  INVX1_477
timestamp 1556798218
transform 1 0 5240 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_415
timestamp 1556798218
transform 1 0 5272 0 1 1810
box 0 0 48 200
use INVX1  INVX1_478
timestamp 1556798218
transform -1 0 5352 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_427
timestamp 1556798218
transform 1 0 5352 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_413
timestamp 1556798218
transform 1 0 5416 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_428
timestamp 1556798218
transform -1 0 5528 0 1 1810
box 0 0 64 200
use INVX1  INVX1_479
timestamp 1556798218
transform -1 0 5560 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_110
timestamp 1556798218
transform 1 0 5560 0 1 1810
box 0 0 64 200
use INVX1  INVX1_438
timestamp 1556798218
transform 1 0 5624 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_394
timestamp 1556798218
transform -1 0 5720 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_259
timestamp 1556798218
transform -1 0 5912 0 1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_260
timestamp 1556798218
transform -1 0 6104 0 1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_150
timestamp 1556798218
transform 1 0 6104 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_228
timestamp 1556798218
transform 1 0 6296 0 1 1810
box 0 0 64 200
use FILL  FILL_9_3_0
timestamp 1556798218
transform -1 0 6376 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_1
timestamp 1556798218
transform -1 0 6392 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_2
timestamp 1556798218
transform -1 0 6408 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_227
timestamp 1556798218
transform -1 0 6472 0 1 1810
box 0 0 64 200
use INVX1  INVX1_244
timestamp 1556798218
transform -1 0 6504 0 1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_75
timestamp 1556798218
transform -1 0 6584 0 1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_92
timestamp 1556798218
transform 1 0 6584 0 1 1810
box 0 0 48 200
use INVX1  INVX1_246
timestamp 1556798218
transform -1 0 6664 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_104
timestamp 1556798218
transform -1 0 6728 0 1 1810
box 0 0 64 200
use INVX1  INVX1_455
timestamp 1556798218
transform 1 0 6728 0 1 1810
box 0 0 32 200
use INVX1  INVX1_457
timestamp 1556798218
transform -1 0 6792 0 1 1810
box 0 0 32 200
use INVX1  INVX1_454
timestamp 1556798218
transform -1 0 6824 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_409
timestamp 1556798218
transform 1 0 6824 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_395
timestamp 1556798218
transform 1 0 6888 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_273
timestamp 1556798218
transform 1 0 6936 0 1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1556798218
transform 1 0 7128 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_33
timestamp 1556798218
transform -1 0 7384 0 1 1810
box 0 0 64 200
use INVX1  INVX1_36
timestamp 1556798218
transform -1 0 7416 0 1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_10
timestamp 1556798218
transform -1 0 7496 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_55
timestamp 1556798218
transform -1 0 7544 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1556798218
transform 1 0 7544 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_39
timestamp 1556798218
transform -1 0 7800 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_57
timestamp 1556798218
transform -1 0 7848 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_41
timestamp 1556798218
transform 1 0 7848 0 1 1810
box 0 0 64 200
use BUFX2  BUFX2_141
timestamp 1556798218
transform 1 0 7912 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_54
timestamp 1556798218
transform -1 0 8008 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_38
timestamp 1556798218
transform 1 0 8008 0 1 1810
box 0 0 64 200
use BUFX2  BUFX2_139
timestamp 1556798218
transform 1 0 8072 0 1 1810
box 0 0 48 200
use FILL  FILL_10_1
timestamp 1556798218
transform 1 0 8120 0 1 1810
box 0 0 16 200
use FILL  FILL_10_2
timestamp 1556798218
transform 1 0 8136 0 1 1810
box 0 0 16 200
use FILL  FILL_10_3
timestamp 1556798218
transform 1 0 8152 0 1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_55
timestamp 1556798218
transform -1 0 72 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_151
timestamp 1556798218
transform 1 0 72 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_161
timestamp 1556798218
transform -1 0 168 0 -1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_65
timestamp 1556798218
transform 1 0 168 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_159
timestamp 1556798218
transform -1 0 248 0 -1 1810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_102
timestamp 1556798218
transform 1 0 248 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_154
timestamp 1556798218
transform -1 0 504 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_164
timestamp 1556798218
transform -1 0 536 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_397
timestamp 1556798218
transform 1 0 536 0 -1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_149
timestamp 1556798218
transform -1 0 616 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_363
timestamp 1556798218
transform -1 0 680 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_353
timestamp 1556798218
transform -1 0 728 0 -1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_58
timestamp 1556798218
transform -1 0 792 0 -1 1810
box 0 0 64 200
use XNOR2X1  XNOR2X1_53
timestamp 1556798218
transform -1 0 904 0 -1 1810
box 0 0 112 200
use INVX1  INVX1_401
timestamp 1556798218
transform -1 0 936 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_398
timestamp 1556798218
transform -1 0 968 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_355
timestamp 1556798218
transform 1 0 968 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_356
timestamp 1556798218
transform -1 0 1064 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_361
timestamp 1556798218
transform 1 0 1064 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_238
timestamp 1556798218
transform -1 0 1320 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_362
timestamp 1556798218
transform -1 0 1384 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_352
timestamp 1556798218
transform -1 0 1432 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_402
timestamp 1556798218
transform -1 0 1464 0 -1 1810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_76
timestamp 1556798218
transform -1 0 1656 0 -1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_140
timestamp 1556798218
transform 1 0 1656 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_113
timestamp 1556798218
transform -1 0 1768 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1556798218
transform -1 0 1784 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1556798218
transform -1 0 1800 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_2
timestamp 1556798218
transform -1 0 1816 0 -1 1810
box 0 0 16 200
use INVX1  INVX1_116
timestamp 1556798218
transform -1 0 1848 0 -1 1810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_75
timestamp 1556798218
transform 1 0 1848 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_101
timestamp 1556798218
transform -1 0 2104 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_114
timestamp 1556798218
transform 1 0 2104 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_115
timestamp 1556798218
transform 1 0 2152 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_79
timestamp 1556798218
transform -1 0 2392 0 -1 1810
box 0 0 192 200
use AOI21X1  AOI21X1_18
timestamp 1556798218
transform -1 0 2456 0 -1 1810
box 0 0 64 200
use XNOR2X1  XNOR2X1_13
timestamp 1556798218
transform 1 0 2456 0 -1 1810
box 0 0 112 200
use NAND3X1  NAND3X1_42
timestamp 1556798218
transform 1 0 2568 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_123
timestamp 1556798218
transform 1 0 2632 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_121
timestamp 1556798218
transform -1 0 2696 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_119
timestamp 1556798218
transform 1 0 2696 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_112
timestamp 1556798218
transform 1 0 2760 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_38
timestamp 1556798218
transform 1 0 2808 0 -1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_128
timestamp 1556798218
transform -1 0 2936 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_116
timestamp 1556798218
transform 1 0 2936 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_117
timestamp 1556798218
transform -1 0 3064 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_53
timestamp 1556798218
transform -1 0 3112 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_39
timestamp 1556798218
transform -1 0 3192 0 -1 1810
box 0 0 80 200
use INVX1  INVX1_122
timestamp 1556798218
transform -1 0 3224 0 -1 1810
box 0 0 32 200
use AND2X2  AND2X2_42
timestamp 1556798218
transform -1 0 3288 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_1_0
timestamp 1556798218
transform 1 0 3288 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1556798218
transform 1 0 3304 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_2
timestamp 1556798218
transform 1 0 3320 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_380
timestamp 1556798218
transform 1 0 3336 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_370
timestamp 1556798218
transform -1 0 3448 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_379
timestamp 1556798218
transform -1 0 3512 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_125
timestamp 1556798218
transform -1 0 3592 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_162
timestamp 1556798218
transform 1 0 3592 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_419
timestamp 1556798218
transform 1 0 3640 0 -1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_124
timestamp 1556798218
transform 1 0 3672 0 -1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_372
timestamp 1556798218
transform 1 0 3752 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_421
timestamp 1556798218
transform -1 0 3832 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_422
timestamp 1556798218
transform -1 0 3864 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_373
timestamp 1556798218
transform 1 0 3864 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_374
timestamp 1556798218
transform -1 0 3960 0 -1 1810
box 0 0 48 200
use BUFX2  BUFX2_28
timestamp 1556798218
transform -1 0 4008 0 -1 1810
box 0 0 48 200
use AND2X2  AND2X2_16
timestamp 1556798218
transform 1 0 4008 0 -1 1810
box 0 0 64 200
use BUFX2  BUFX2_111
timestamp 1556798218
transform 1 0 4072 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_335
timestamp 1556798218
transform -1 0 4312 0 -1 1810
box 0 0 192 200
use INVX1  INVX1_571
timestamp 1556798218
transform 1 0 4312 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_508
timestamp 1556798218
transform 1 0 4344 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_418
timestamp 1556798218
transform -1 0 4472 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_337
timestamp 1556798218
transform 1 0 4472 0 -1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_177
timestamp 1556798218
transform -1 0 4712 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_275
timestamp 1556798218
transform -1 0 4904 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_2_0
timestamp 1556798218
transform 1 0 4904 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1556798218
transform 1 0 4920 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_2
timestamp 1556798218
transform 1 0 4936 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_400
timestamp 1556798218
transform 1 0 4952 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_402
timestamp 1556798218
transform 1 0 5000 0 -1 1810
box 0 0 48 200
use NOR3X1  NOR3X1_5
timestamp 1556798218
transform 1 0 5048 0 -1 1810
box 0 0 128 200
use NAND2X1  NAND2X1_401
timestamp 1556798218
transform 1 0 5176 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_414
timestamp 1556798218
transform -1 0 5272 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_140
timestamp 1556798218
transform -1 0 5352 0 -1 1810
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_284
timestamp 1556798218
transform 1 0 5352 0 -1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_417
timestamp 1556798218
transform 1 0 5544 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_416
timestamp 1556798218
transform -1 0 5640 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_141
timestamp 1556798218
transform 1 0 5640 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_184
timestamp 1556798218
transform -1 0 5768 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_282
timestamp 1556798218
transform 1 0 5768 0 -1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_87
timestamp 1556798218
transform 1 0 5960 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_229
timestamp 1556798218
transform -1 0 6040 0 -1 1810
box 0 0 32 200
use BUFX2  BUFX2_34
timestamp 1556798218
transform -1 0 6088 0 -1 1810
box 0 0 48 200
use BUFX2  BUFX2_31
timestamp 1556798218
transform 1 0 6088 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_153
timestamp 1556798218
transform -1 0 6328 0 -1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_228
timestamp 1556798218
transform -1 0 6376 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_3_0
timestamp 1556798218
transform -1 0 6392 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_1
timestamp 1556798218
transform -1 0 6408 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_2
timestamp 1556798218
transform -1 0 6424 0 -1 1810
box 0 0 16 200
use INVX1  INVX1_245
timestamp 1556798218
transform -1 0 6456 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_225
timestamp 1556798218
transform -1 0 6520 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_74
timestamp 1556798218
transform 1 0 6520 0 -1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_78
timestamp 1556798218
transform 1 0 6600 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_230
timestamp 1556798218
transform 1 0 6664 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_247
timestamp 1556798218
transform -1 0 6744 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_231
timestamp 1556798218
transform 1 0 6744 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_232
timestamp 1556798218
transform -1 0 6840 0 -1 1810
box 0 0 48 200
use BUFX2  BUFX2_112
timestamp 1556798218
transform -1 0 6888 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_458
timestamp 1556798218
transform 1 0 6888 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_410
timestamp 1556798218
transform 1 0 6920 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_270
timestamp 1556798218
transform -1 0 7176 0 -1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_369
timestamp 1556798218
transform 1 0 7176 0 -1 1810
box 0 0 48 200
use BUFX2  BUFX2_114
timestamp 1556798218
transform 1 0 7224 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_47
timestamp 1556798218
transform 1 0 7272 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_30
timestamp 1556798218
transform -1 0 7384 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1556798218
transform 1 0 7384 0 -1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_269
timestamp 1556798218
transform -1 0 7768 0 -1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1556798218
transform 1 0 7768 0 -1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1556798218
transform 1 0 7960 0 -1 1810
box 0 0 192 200
use FILL  FILL_9_1
timestamp 1556798218
transform -1 0 8168 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_54
timestamp 1556798218
transform -1 0 72 0 1 1410
box 0 0 64 200
use INVX1  INVX1_162
timestamp 1556798218
transform 1 0 72 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_152
timestamp 1556798218
transform -1 0 168 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_155
timestamp 1556798218
transform -1 0 232 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_161
timestamp 1556798218
transform -1 0 280 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_66
timestamp 1556798218
transform 1 0 280 0 1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_50
timestamp 1556798218
transform -1 0 408 0 1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_153
timestamp 1556798218
transform 1 0 408 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_51
timestamp 1556798218
transform -1 0 552 0 1 1410
box 0 0 80 200
use INVX1  INVX1_160
timestamp 1556798218
transform -1 0 584 0 1 1410
box 0 0 32 200
use AND2X2  AND2X2_49
timestamp 1556798218
transform -1 0 648 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_94
timestamp 1556798218
transform -1 0 712 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_240
timestamp 1556798218
transform 1 0 712 0 1 1410
box 0 0 192 200
use BUFX2  BUFX2_41
timestamp 1556798218
transform 1 0 904 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_74
timestamp 1556798218
transform 1 0 952 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_111
timestamp 1556798218
transform 1 0 1144 0 1 1410
box 0 0 64 200
use INVX1  INVX1_115
timestamp 1556798218
transform -1 0 1240 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_110
timestamp 1556798218
transform -1 0 1304 0 1 1410
box 0 0 64 200
use INVX1  INVX1_114
timestamp 1556798218
transform 1 0 1304 0 1 1410
box 0 0 32 200
use AND2X2  AND2X2_41
timestamp 1556798218
transform 1 0 1336 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_37
timestamp 1556798218
transform 1 0 1400 0 1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_51
timestamp 1556798218
transform 1 0 1480 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_40
timestamp 1556798218
transform -1 0 1592 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_122
timestamp 1556798218
transform 1 0 1592 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_17
timestamp 1556798218
transform -1 0 1704 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_36
timestamp 1556798218
transform 1 0 1704 0 1 1410
box 0 0 80 200
use FILL  FILL_7_0_0
timestamp 1556798218
transform -1 0 1800 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1556798218
transform -1 0 1816 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_2
timestamp 1556798218
transform -1 0 1832 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_123
timestamp 1556798218
transform -1 0 1880 0 1 1410
box 0 0 48 200
use INVX1  INVX1_113
timestamp 1556798218
transform -1 0 1912 0 1 1410
box 0 0 32 200
use XNOR2X1  XNOR2X1_12
timestamp 1556798218
transform -1 0 2024 0 1 1410
box 0 0 112 200
use INVX1  INVX1_416
timestamp 1556798218
transform -1 0 2056 0 1 1410
box 0 0 32 200
use AND2X2  AND2X2_95
timestamp 1556798218
transform 1 0 2056 0 1 1410
box 0 0 64 200
use BUFX2  BUFX2_103
timestamp 1556798218
transform -1 0 2168 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_366
timestamp 1556798218
transform 1 0 2168 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_365
timestamp 1556798218
transform 1 0 2216 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_41
timestamp 1556798218
transform 1 0 2264 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_106
timestamp 1556798218
transform 1 0 2312 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_80
timestamp 1556798218
transform 1 0 2360 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_98
timestamp 1556798218
transform -1 0 2600 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_78
timestamp 1556798218
transform 1 0 2600 0 1 1410
box 0 0 192 200
use BUFX2  BUFX2_72
timestamp 1556798218
transform -1 0 2840 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_252
timestamp 1556798218
transform 1 0 2840 0 1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_250
timestamp 1556798218
transform 1 0 3032 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_382
timestamp 1556798218
transform -1 0 3288 0 1 1410
box 0 0 64 200
use FILL  FILL_7_1_0
timestamp 1556798218
transform -1 0 3304 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1556798218
transform -1 0 3320 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_2
timestamp 1556798218
transform -1 0 3336 0 1 1410
box 0 0 16 200
use INVX1  INVX1_424
timestamp 1556798218
transform -1 0 3368 0 1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_251
timestamp 1556798218
transform 1 0 3368 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_368
timestamp 1556798218
transform 1 0 3560 0 1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_4
timestamp 1556798218
transform -1 0 3736 0 1 1410
box 0 0 128 200
use NAND2X1  NAND2X1_367
timestamp 1556798218
transform -1 0 3784 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_179
timestamp 1556798218
transform 1 0 3784 0 1 1410
box 0 0 48 200
use INVX1  INVX1_460
timestamp 1556798218
transform -1 0 3864 0 1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_274
timestamp 1556798218
transform 1 0 3864 0 1 1410
box 0 0 192 200
use AOI22X1  AOI22X1_137
timestamp 1556798218
transform -1 0 4136 0 1 1410
box 0 0 80 200
use NAND2X1  NAND2X1_407
timestamp 1556798218
transform -1 0 4184 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_416
timestamp 1556798218
transform 1 0 4184 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_415
timestamp 1556798218
transform -1 0 4312 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_403
timestamp 1556798218
transform -1 0 4360 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_405
timestamp 1556798218
transform -1 0 4408 0 1 1410
box 0 0 48 200
use INVX1  INVX1_464
timestamp 1556798218
transform -1 0 4440 0 1 1410
box 0 0 32 200
use INVX1  INVX1_461
timestamp 1556798218
transform 1 0 4440 0 1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_276
timestamp 1556798218
transform 1 0 4472 0 1 1410
box 0 0 192 200
use AND2X2  AND2X2_106
timestamp 1556798218
transform -1 0 4728 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_175
timestamp 1556798218
transform -1 0 4776 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_133
timestamp 1556798218
transform -1 0 4824 0 1 1410
box 0 0 48 200
use FILL  FILL_7_2_0
timestamp 1556798218
transform 1 0 4824 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1556798218
transform 1 0 4840 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_2
timestamp 1556798218
transform 1 0 4856 0 1 1410
box 0 0 16 200
use AND2X2  AND2X2_105
timestamp 1556798218
transform 1 0 4872 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_173
timestamp 1556798218
transform -1 0 4984 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_283
timestamp 1556798218
transform -1 0 5176 0 1 1410
box 0 0 192 200
use INVX1  INVX1_480
timestamp 1556798218
transform 1 0 5176 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_430
timestamp 1556798218
transform 1 0 5208 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_145
timestamp 1556798218
transform -1 0 5464 0 1 1410
box 0 0 192 200
use AND2X2  AND2X2_97
timestamp 1556798218
transform 1 0 5464 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_158
timestamp 1556798218
transform -1 0 5576 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_219
timestamp 1556798218
transform 1 0 5576 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_217
timestamp 1556798218
transform 1 0 5624 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_75
timestamp 1556798218
transform 1 0 5688 0 1 1410
box 0 0 64 200
use INVX1  INVX1_231
timestamp 1556798218
transform -1 0 5784 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_213
timestamp 1556798218
transform -1 0 5848 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_214
timestamp 1556798218
transform -1 0 5912 0 1 1410
box 0 0 64 200
use CLKBUF1  CLKBUF1_35
timestamp 1556798218
transform -1 0 6056 0 1 1410
box 0 0 144 200
use BUFX2  BUFX2_5
timestamp 1556798218
transform -1 0 6104 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_226
timestamp 1556798218
transform 1 0 6104 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_36
timestamp 1556798218
transform 1 0 6168 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_79
timestamp 1556798218
transform -1 0 6296 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_229
timestamp 1556798218
transform -1 0 6360 0 1 1410
box 0 0 64 200
use FILL  FILL_7_3_0
timestamp 1556798218
transform -1 0 6376 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_1
timestamp 1556798218
transform -1 0 6392 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_2
timestamp 1556798218
transform -1 0 6408 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_229
timestamp 1556798218
transform -1 0 6456 0 1 1410
box 0 0 48 200
use INVX1  INVX1_249
timestamp 1556798218
transform 1 0 6456 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_230
timestamp 1556798218
transform 1 0 6488 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_151
timestamp 1556798218
transform -1 0 6744 0 1 1410
box 0 0 192 200
use INVX1  INVX1_225
timestamp 1556798218
transform 1 0 6744 0 1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_214
timestamp 1556798218
transform -1 0 6824 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_215
timestamp 1556798218
transform -1 0 6872 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_86
timestamp 1556798218
transform -1 0 6920 0 1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_69
timestamp 1556798218
transform -1 0 7000 0 1 1410
box 0 0 80 200
use INVX1  INVX1_228
timestamp 1556798218
transform 1 0 7000 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_211
timestamp 1556798218
transform 1 0 7032 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_139
timestamp 1556798218
transform -1 0 7288 0 1 1410
box 0 0 192 200
use CLKBUF1  CLKBUF1_6
timestamp 1556798218
transform 1 0 7288 0 1 1410
box 0 0 144 200
use BUFX2  BUFX2_113
timestamp 1556798218
transform 1 0 7432 0 1 1410
box 0 0 48 200
use AND2X2  AND2X2_103
timestamp 1556798218
transform 1 0 7480 0 1 1410
box 0 0 64 200
use INVX1  INVX1_451
timestamp 1556798218
transform 1 0 7544 0 1 1410
box 0 0 32 200
use INVX1  INVX1_446
timestamp 1556798218
transform 1 0 7576 0 1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_169
timestamp 1556798218
transform -1 0 7656 0 1 1410
box 0 0 48 200
use INVX1  INVX1_447
timestamp 1556798218
transform 1 0 7656 0 1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_137
timestamp 1556798218
transform 1 0 7688 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_402
timestamp 1556798218
transform 1 0 7752 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_405
timestamp 1556798218
transform -1 0 7880 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_401
timestamp 1556798218
transform 1 0 7880 0 1 1410
box 0 0 64 200
use INVX1  INVX1_449
timestamp 1556798218
transform -1 0 7976 0 1 1410
box 0 0 32 200
use INVX1  INVX1_448
timestamp 1556798218
transform -1 0 8008 0 1 1410
box 0 0 32 200
use XNOR2X1  XNOR2X1_60
timestamp 1556798218
transform -1 0 8120 0 1 1410
box 0 0 112 200
use FILL  FILL_8_1
timestamp 1556798218
transform 1 0 8120 0 1 1410
box 0 0 16 200
use FILL  FILL_8_2
timestamp 1556798218
transform 1 0 8136 0 1 1410
box 0 0 16 200
use FILL  FILL_8_3
timestamp 1556798218
transform 1 0 8152 0 1 1410
box 0 0 16 200
use XNOR2X1  XNOR2X1_19
timestamp 1556798218
transform -1 0 120 0 -1 1410
box 0 0 112 200
use AOI21X1  AOI21X1_24
timestamp 1556798218
transform 1 0 120 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_104
timestamp 1556798218
transform 1 0 184 0 -1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_162
timestamp 1556798218
transform -1 0 424 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_163
timestamp 1556798218
transform -1 0 456 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_163
timestamp 1556798218
transform 1 0 456 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_164
timestamp 1556798218
transform -1 0 552 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_160
timestamp 1556798218
transform -1 0 600 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_362
timestamp 1556798218
transform 1 0 600 0 -1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_133
timestamp 1556798218
transform -1 0 680 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_221
timestamp 1556798218
transform 1 0 680 0 -1 1410
box 0 0 192 200
use CLKBUF1  CLKBUF1_30
timestamp 1556798218
transform -1 0 1016 0 -1 1410
box 0 0 144 200
use NAND2X1  NAND2X1_121
timestamp 1556798218
transform 1 0 1016 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_367
timestamp 1556798218
transform -1 0 1096 0 -1 1410
box 0 0 32 200
use AND2X2  AND2X2_4
timestamp 1556798218
transform -1 0 1160 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_111
timestamp 1556798218
transform 1 0 1160 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_124
timestamp 1556798218
transform 1 0 1192 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_125
timestamp 1556798218
transform -1 0 1288 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_336
timestamp 1556798218
transform -1 0 1336 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_112
timestamp 1556798218
transform 1 0 1336 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_108
timestamp 1556798218
transform -1 0 1432 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_109
timestamp 1556798218
transform -1 0 1496 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_97
timestamp 1556798218
transform 1 0 1496 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_41
timestamp 1556798218
transform -1 0 1608 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_112
timestamp 1556798218
transform 1 0 1608 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_0_0
timestamp 1556798218
transform -1 0 1688 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1556798218
transform -1 0 1704 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_2
timestamp 1556798218
transform -1 0 1720 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_246
timestamp 1556798218
transform -1 0 1912 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_374
timestamp 1556798218
transform -1 0 1976 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_373
timestamp 1556798218
transform -1 0 2040 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_415
timestamp 1556798218
transform -1 0 2072 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_362
timestamp 1556798218
transform -1 0 2120 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_303
timestamp 1556798218
transform -1 0 2168 0 -1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_123
timestamp 1556798218
transform 1 0 2168 0 -1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_154
timestamp 1556798218
transform 1 0 2248 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_414
timestamp 1556798218
transform 1 0 2296 0 -1 1410
box 0 0 32 200
use INVX1  INVX1_413
timestamp 1556798218
transform 1 0 2328 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_364
timestamp 1556798218
transform 1 0 2360 0 -1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_122
timestamp 1556798218
transform -1 0 2488 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_249
timestamp 1556798218
transform -1 0 2680 0 -1 1410
box 0 0 192 200
use BUFX2  BUFX2_1
timestamp 1556798218
transform 1 0 2680 0 -1 1410
box 0 0 48 200
use CLKBUF1  CLKBUF1_8
timestamp 1556798218
transform 1 0 2728 0 -1 1410
box 0 0 144 200
use INVX1  INVX1_354
timestamp 1556798218
transform 1 0 2872 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_211
timestamp 1556798218
transform -1 0 3096 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_322
timestamp 1556798218
transform 1 0 3096 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_210
timestamp 1556798218
transform 1 0 3160 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_1_0
timestamp 1556798218
transform -1 0 3368 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1556798218
transform -1 0 3384 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_2
timestamp 1556798218
transform -1 0 3400 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_320
timestamp 1556798218
transform -1 0 3464 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_314
timestamp 1556798218
transform -1 0 3512 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_353
timestamp 1556798218
transform -1 0 3544 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_255
timestamp 1556798218
transform 1 0 3544 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_388
timestamp 1556798218
transform -1 0 3800 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_431
timestamp 1556798218
transform -1 0 3832 0 -1 1410
box 0 0 32 200
use AND2X2  AND2X2_108
timestamp 1556798218
transform -1 0 3896 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_465
timestamp 1556798218
transform 1 0 3896 0 -1 1410
box 0 0 32 200
use INVX1  INVX1_463
timestamp 1556798218
transform 1 0 3928 0 -1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_180
timestamp 1556798218
transform -1 0 4008 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_406
timestamp 1556798218
transform 1 0 4008 0 -1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_136
timestamp 1556798218
transform -1 0 4136 0 -1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_140
timestamp 1556798218
transform -1 0 4200 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_141
timestamp 1556798218
transform 1 0 4200 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_414
timestamp 1556798218
transform 1 0 4264 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_413
timestamp 1556798218
transform 1 0 4328 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_67
timestamp 1556798218
transform 1 0 4392 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_417
timestamp 1556798218
transform -1 0 4520 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_404
timestamp 1556798218
transform -1 0 4568 0 -1 1410
box 0 0 48 200
use BUFX2  BUFX2_131
timestamp 1556798218
transform -1 0 4616 0 -1 1410
box 0 0 48 200
use XNOR2X1  XNOR2X1_66
timestamp 1556798218
transform 1 0 4616 0 -1 1410
box 0 0 112 200
use NOR2X1  NOR2X1_176
timestamp 1556798218
transform -1 0 4776 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_492
timestamp 1556798218
transform 1 0 4776 0 -1 1410
box 0 0 32 200
use FILL  FILL_6_2_0
timestamp 1556798218
transform 1 0 4808 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1556798218
transform 1 0 4824 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_2
timestamp 1556798218
transform 1 0 4840 0 -1 1410
box 0 0 16 200
use AOI21X1  AOI21X1_71
timestamp 1556798218
transform 1 0 4856 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_174
timestamp 1556798218
transform -1 0 4968 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_292
timestamp 1556798218
transform 1 0 4968 0 -1 1410
box 0 0 192 200
use NOR2X1  NOR2X1_156
timestamp 1556798218
transform -1 0 5208 0 -1 1410
box 0 0 48 200
use AND2X2  AND2X2_96
timestamp 1556798218
transform -1 0 5272 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_155
timestamp 1556798218
transform -1 0 5320 0 -1 1410
box 0 0 48 200
use XNOR2X1  XNOR2X1_29
timestamp 1556798218
transform -1 0 5432 0 -1 1410
box 0 0 112 200
use AOI21X1  AOI21X1_34
timestamp 1556798218
transform 1 0 5432 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_221
timestamp 1556798218
transform 1 0 5496 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_157
timestamp 1556798218
transform 1 0 5544 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_230
timestamp 1556798218
transform -1 0 5624 0 -1 1410
box 0 0 32 200
use INVX1  INVX1_232
timestamp 1556798218
transform 1 0 5624 0 -1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_74
timestamp 1556798218
transform -1 0 5720 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_159
timestamp 1556798218
transform 1 0 5720 0 -1 1410
box 0 0 48 200
use AND2X2  AND2X2_98
timestamp 1556798218
transform 1 0 5768 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_160
timestamp 1556798218
transform -1 0 5880 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_243
timestamp 1556798218
transform 1 0 5880 0 -1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_91
timestamp 1556798218
transform -1 0 5960 0 -1 1410
box 0 0 48 200
use BUFX2  BUFX2_14
timestamp 1556798218
transform -1 0 6008 0 -1 1410
box 0 0 48 200
use BUFX2  BUFX2_15
timestamp 1556798218
transform 1 0 6008 0 -1 1410
box 0 0 48 200
use XNOR2X1  XNOR2X1_31
timestamp 1556798218
transform 1 0 6056 0 -1 1410
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_152
timestamp 1556798218
transform 1 0 6168 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_3_0
timestamp 1556798218
transform 1 0 6360 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_1
timestamp 1556798218
transform 1 0 6376 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_2
timestamp 1556798218
transform 1 0 6392 0 -1 1410
box 0 0 16 200
use BUFX2  BUFX2_67
timestamp 1556798218
transform 1 0 6408 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_206
timestamp 1556798218
transform 1 0 6456 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_207
timestamp 1556798218
transform -1 0 6584 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_213
timestamp 1556798218
transform 1 0 6584 0 -1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_68
timestamp 1556798218
transform -1 0 6712 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_138
timestamp 1556798218
transform 1 0 6712 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_208
timestamp 1556798218
transform 1 0 6904 0 -1 1410
box 0 0 64 200
use CLKBUF1  CLKBUF1_45
timestamp 1556798218
transform 1 0 6968 0 -1 1410
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_115
timestamp 1556798218
transform -1 0 7304 0 -1 1410
box 0 0 192 200
use INVX1  INVX1_186
timestamp 1556798218
transform 1 0 7304 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_266
timestamp 1556798218
transform 1 0 7336 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_404
timestamp 1556798218
transform -1 0 7592 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_390
timestamp 1556798218
transform 1 0 7592 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_403
timestamp 1556798218
transform -1 0 7704 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_450
timestamp 1556798218
transform 1 0 7704 0 -1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_136
timestamp 1556798218
transform 1 0 7736 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_391
timestamp 1556798218
transform 1 0 7800 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_392
timestamp 1556798218
transform 1 0 7848 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_65
timestamp 1556798218
transform -1 0 7960 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_268
timestamp 1556798218
transform 1 0 7960 0 -1 1410
box 0 0 192 200
use FILL  FILL_7_1
timestamp 1556798218
transform -1 0 8168 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_244
timestamp 1556798218
transform -1 0 200 0 1 1010
box 0 0 192 200
use XNOR2X1  XNOR2X1_54
timestamp 1556798218
transform -1 0 312 0 1 1010
box 0 0 112 200
use BUFX2  BUFX2_39
timestamp 1556798218
transform -1 0 360 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_48
timestamp 1556798218
transform -1 0 408 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_156
timestamp 1556798218
transform 1 0 408 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_220
timestamp 1556798218
transform 1 0 472 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_333
timestamp 1556798218
transform -1 0 728 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_113
timestamp 1556798218
transform 1 0 728 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_325
timestamp 1556798218
transform 1 0 792 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_330
timestamp 1556798218
transform 1 0 840 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_329
timestamp 1556798218
transform -1 0 968 0 1 1010
box 0 0 64 200
use INVX1  INVX1_363
timestamp 1556798218
transform -1 0 1000 0 1 1010
box 0 0 32 200
use INVX1  INVX1_364
timestamp 1556798218
transform -1 0 1032 0 1 1010
box 0 0 32 200
use INVX1  INVX1_365
timestamp 1556798218
transform 1 0 1032 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_134
timestamp 1556798218
transform -1 0 1112 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_109
timestamp 1556798218
transform -1 0 1192 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_328
timestamp 1556798218
transform 1 0 1192 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_327
timestamp 1556798218
transform -1 0 1288 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_119
timestamp 1556798218
transform -1 0 1336 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_2
timestamp 1556798218
transform 1 0 1336 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_117
timestamp 1556798218
transform 1 0 1400 0 1 1010
box 0 0 48 200
use INVX1  INVX1_106
timestamp 1556798218
transform 1 0 1448 0 1 1010
box 0 0 32 200
use INVX1  INVX1_104
timestamp 1556798218
transform -1 0 1512 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_116
timestamp 1556798218
transform 1 0 1512 0 1 1010
box 0 0 48 200
use XNOR2X1  XNOR2X1_11
timestamp 1556798218
transform -1 0 1672 0 1 1010
box 0 0 112 200
use NAND2X1  NAND2X1_119
timestamp 1556798218
transform 1 0 1672 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_120
timestamp 1556798218
transform -1 0 1768 0 1 1010
box 0 0 48 200
use FILL  FILL_5_0_0
timestamp 1556798218
transform -1 0 1784 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1556798218
transform -1 0 1800 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_2
timestamp 1556798218
transform -1 0 1816 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_77
timestamp 1556798218
transform -1 0 2008 0 1 1010
box 0 0 192 200
use INVX1  INVX1_110
timestamp 1556798218
transform 1 0 2008 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_50
timestamp 1556798218
transform -1 0 2088 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_40
timestamp 1556798218
transform 1 0 2088 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_60
timestamp 1556798218
transform 1 0 2136 0 1 1010
box 0 0 64 200
use XNOR2X1  XNOR2X1_55
timestamp 1556798218
transform -1 0 2312 0 1 1010
box 0 0 112 200
use INVX1  INVX1_412
timestamp 1556798218
transform -1 0 2344 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_375
timestamp 1556798218
transform 1 0 2344 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_363
timestamp 1556798218
transform -1 0 2456 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_126
timestamp 1556798218
transform -1 0 2520 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_371
timestamp 1556798218
transform 1 0 2520 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_372
timestamp 1556798218
transform -1 0 2648 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_127
timestamp 1556798218
transform 1 0 2648 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_153
timestamp 1556798218
transform 1 0 2712 0 1 1010
box 0 0 48 200
use INVX1  INVX1_411
timestamp 1556798218
transform -1 0 2792 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_376
timestamp 1556798218
transform -1 0 2856 0 1 1010
box 0 0 64 200
use INVX1  INVX1_417
timestamp 1556798218
transform -1 0 2888 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_247
timestamp 1556798218
transform 1 0 2888 0 1 1010
box 0 0 192 200
use CLKBUF1  CLKBUF1_36
timestamp 1556798218
transform 1 0 3080 0 1 1010
box 0 0 144 200
use AOI22X1  AOI22X1_104
timestamp 1556798218
transform 1 0 3224 0 1 1010
box 0 0 80 200
use FILL  FILL_5_1_0
timestamp 1556798218
transform 1 0 3304 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1556798218
transform 1 0 3320 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_2
timestamp 1556798218
transform 1 0 3336 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_316
timestamp 1556798218
transform 1 0 3352 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_319
timestamp 1556798218
transform -1 0 3464 0 1 1010
box 0 0 64 200
use INVX1  INVX1_349
timestamp 1556798218
transform 1 0 3464 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_130
timestamp 1556798218
transform -1 0 3544 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_105
timestamp 1556798218
transform -1 0 3624 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_318
timestamp 1556798218
transform -1 0 3672 0 1 1010
box 0 0 48 200
use INVX1  INVX1_352
timestamp 1556798218
transform -1 0 3704 0 1 1010
box 0 0 32 200
use AND2X2  AND2X2_83
timestamp 1556798218
transform 1 0 3704 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_212
timestamp 1556798218
transform -1 0 3960 0 1 1010
box 0 0 192 200
use AOI22X1  AOI22X1_127
timestamp 1556798218
transform -1 0 4040 0 1 1010
box 0 0 80 200
use AND2X2  AND2X2_100
timestamp 1556798218
transform -1 0 4104 0 1 1010
box 0 0 64 200
use INVX1  INVX1_426
timestamp 1556798218
transform 1 0 4104 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_164
timestamp 1556798218
transform 1 0 4136 0 1 1010
box 0 0 48 200
use INVX1  INVX1_428
timestamp 1556798218
transform -1 0 4216 0 1 1010
box 0 0 32 200
use AOI22X1  AOI22X1_126
timestamp 1556798218
transform -1 0 4296 0 1 1010
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_277
timestamp 1556798218
transform 1 0 4296 0 1 1010
box 0 0 192 200
use INVX1  INVX1_462
timestamp 1556798218
transform -1 0 4520 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_290
timestamp 1556798218
transform -1 0 4712 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_440
timestamp 1556798218
transform 1 0 4712 0 1 1010
box 0 0 64 200
use INVX1  INVX1_493
timestamp 1556798218
transform -1 0 4808 0 1 1010
box 0 0 32 200
use FILL  FILL_5_2_0
timestamp 1556798218
transform -1 0 4824 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1556798218
transform -1 0 4840 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_2
timestamp 1556798218
transform -1 0 4856 0 1 1010
box 0 0 16 200
use AND2X2  AND2X2_112
timestamp 1556798218
transform -1 0 4920 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_439
timestamp 1556798218
transform -1 0 4984 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_425
timestamp 1556798218
transform -1 0 5032 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_148
timestamp 1556798218
transform -1 0 5096 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_437
timestamp 1556798218
transform 1 0 5096 0 1 1010
box 0 0 64 200
use INVX1  INVX1_490
timestamp 1556798218
transform -1 0 5192 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_441
timestamp 1556798218
transform 1 0 5192 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_424
timestamp 1556798218
transform -1 0 5304 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_438
timestamp 1556798218
transform -1 0 5368 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_149
timestamp 1556798218
transform 1 0 5368 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_293
timestamp 1556798218
transform -1 0 5624 0 1 1010
box 0 0 192 200
use INVX1  INVX1_234
timestamp 1556798218
transform 1 0 5624 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_216
timestamp 1556798218
transform 1 0 5656 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_218
timestamp 1556798218
transform -1 0 5768 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_215
timestamp 1556798218
transform -1 0 5832 0 1 1010
box 0 0 64 200
use INVX1  INVX1_233
timestamp 1556798218
transform -1 0 5864 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_222
timestamp 1556798218
transform 1 0 5864 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_220
timestamp 1556798218
transform -1 0 5960 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_61
timestamp 1556798218
transform 1 0 5960 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_71
timestamp 1556798218
transform 1 0 6024 0 1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_88
timestamp 1556798218
transform 1 0 6104 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_70
timestamp 1556798218
transform -1 0 6232 0 1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_218
timestamp 1556798218
transform -1 0 6296 0 1 1010
box 0 0 64 200
use INVX1  INVX1_235
timestamp 1556798218
transform -1 0 6328 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_80
timestamp 1556798218
transform 1 0 6328 0 1 1010
box 0 0 48 200
use FILL  FILL_5_3_0
timestamp 1556798218
transform 1 0 6376 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_1
timestamp 1556798218
transform 1 0 6392 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_2
timestamp 1556798218
transform 1 0 6408 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_143
timestamp 1556798218
transform 1 0 6424 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_200
timestamp 1556798218
transform -1 0 6664 0 1 1010
box 0 0 48 200
use INVX1  INVX1_224
timestamp 1556798218
transform 1 0 6664 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_212
timestamp 1556798218
transform -1 0 6744 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_73
timestamp 1556798218
transform 1 0 6744 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_72
timestamp 1556798218
transform 1 0 6808 0 1 1010
box 0 0 64 200
use INVX1  INVX1_223
timestamp 1556798218
transform 1 0 6872 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_141
timestamp 1556798218
transform 1 0 6904 0 1 1010
box 0 0 192 200
use AND2X2  AND2X2_60
timestamp 1556798218
transform -1 0 7160 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_211
timestamp 1556798218
transform 1 0 7160 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_209
timestamp 1556798218
transform -1 0 7272 0 1 1010
box 0 0 64 200
use INVX1  INVX1_227
timestamp 1556798218
transform 1 0 7272 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_174
timestamp 1556798218
transform -1 0 7368 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_180
timestamp 1556798218
transform -1 0 7416 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_56
timestamp 1556798218
transform 1 0 7416 0 1 1010
box 0 0 80 200
use INVX1  INVX1_182
timestamp 1556798218
transform 1 0 7496 0 1 1010
box 0 0 32 200
use INVX1  INVX1_183
timestamp 1556798218
transform -1 0 7560 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_169
timestamp 1556798218
transform 1 0 7560 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_170
timestamp 1556798218
transform -1 0 7688 0 1 1010
box 0 0 64 200
use INVX1  INVX1_181
timestamp 1556798218
transform -1 0 7720 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_178
timestamp 1556798218
transform -1 0 7768 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_72
timestamp 1556798218
transform 1 0 7768 0 1 1010
box 0 0 48 200
use INVX1  INVX1_180
timestamp 1556798218
transform 1 0 7816 0 1 1010
box 0 0 32 200
use AOI22X1  AOI22X1_132
timestamp 1556798218
transform 1 0 7848 0 1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_170
timestamp 1556798218
transform -1 0 7976 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_133
timestamp 1556798218
transform -1 0 8056 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_394
timestamp 1556798218
transform 1 0 8056 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_393
timestamp 1556798218
transform 1 0 8104 0 1 1010
box 0 0 48 200
use FILL  FILL_6_1
timestamp 1556798218
transform 1 0 8152 0 1 1010
box 0 0 16 200
use INVX1  INVX1_408
timestamp 1556798218
transform 1 0 8 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_358
timestamp 1556798218
transform 1 0 40 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_59
timestamp 1556798218
transform 1 0 88 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_369
timestamp 1556798218
transform 1 0 152 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_406
timestamp 1556798218
transform -1 0 248 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_365
timestamp 1556798218
transform -1 0 312 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_366
timestamp 1556798218
transform -1 0 376 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_125
timestamp 1556798218
transform -1 0 440 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_151
timestamp 1556798218
transform 1 0 440 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_404
timestamp 1556798218
transform -1 0 520 0 -1 1010
box 0 0 32 200
use INVX1  INVX1_409
timestamp 1556798218
transform -1 0 552 0 -1 1010
box 0 0 32 200
use AOI21X1  AOI21X1_53
timestamp 1556798218
transform -1 0 616 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_366
timestamp 1556798218
transform -1 0 648 0 -1 1010
box 0 0 32 200
use XNOR2X1  XNOR2X1_48
timestamp 1556798218
transform 1 0 648 0 -1 1010
box 0 0 112 200
use NAND3X1  NAND3X1_112
timestamp 1556798218
transform 1 0 760 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_326
timestamp 1556798218
transform 1 0 824 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_108
timestamp 1556798218
transform -1 0 952 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_331
timestamp 1556798218
transform 1 0 952 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_332
timestamp 1556798218
transform -1 0 1080 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_324
timestamp 1556798218
transform -1 0 1128 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_334
timestamp 1556798218
transform -1 0 1192 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_105
timestamp 1556798218
transform -1 0 1224 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_102
timestamp 1556798218
transform -1 0 1288 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_106
timestamp 1556798218
transform 1 0 1288 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_103
timestamp 1556798218
transform -1 0 1416 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1556798218
transform 1 0 1416 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_104
timestamp 1556798218
transform 1 0 1480 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_16
timestamp 1556798218
transform -1 0 1608 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_118
timestamp 1556798218
transform 1 0 1608 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_34
timestamp 1556798218
transform -1 0 1736 0 -1 1010
box 0 0 80 200
use FILL  FILL_4_0_0
timestamp 1556798218
transform -1 0 1752 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1556798218
transform -1 0 1768 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_2
timestamp 1556798218
transform -1 0 1784 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_107
timestamp 1556798218
transform -1 0 1816 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_72
timestamp 1556798218
transform -1 0 2008 0 -1 1010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_248
timestamp 1556798218
transform -1 0 2200 0 -1 1010
box 0 0 192 200
use AND2X2  AND2X2_6
timestamp 1556798218
transform 1 0 2200 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_93
timestamp 1556798218
transform -1 0 2456 0 -1 1010
box 0 0 192 200
use NOR2X1  NOR2X1_59
timestamp 1556798218
transform 1 0 2456 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_138
timestamp 1556798218
transform -1 0 2536 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_146
timestamp 1556798218
transform 1 0 2536 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_147
timestamp 1556798218
transform -1 0 2632 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_137
timestamp 1556798218
transform 1 0 2632 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_144
timestamp 1556798218
transform -1 0 2728 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_91
timestamp 1556798218
transform 1 0 2728 0 -1 1010
box 0 0 192 200
use INVX1  INVX1_351
timestamp 1556798218
transform 1 0 2920 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_317
timestamp 1556798218
transform 1 0 2952 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_318
timestamp 1556798218
transform -1 0 3080 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_315
timestamp 1556798218
transform 1 0 3080 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_321
timestamp 1556798218
transform 1 0 3128 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_350
timestamp 1556798218
transform -1 0 3224 0 -1 1010
box 0 0 32 200
use AOI21X1  AOI21X1_51
timestamp 1556798218
transform -1 0 3288 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_1_0
timestamp 1556798218
transform 1 0 3288 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1556798218
transform 1 0 3304 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_2
timestamp 1556798218
transform 1 0 3320 0 -1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_108
timestamp 1556798218
transform 1 0 3336 0 -1 1010
box 0 0 64 200
use XNOR2X1  XNOR2X1_46
timestamp 1556798218
transform 1 0 3400 0 -1 1010
box 0 0 112 200
use BUFX2  BUFX2_84
timestamp 1556798218
transform -1 0 3560 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_86
timestamp 1556798218
transform -1 0 3608 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_317
timestamp 1556798218
transform 1 0 3608 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_87
timestamp 1556798218
transform 1 0 3656 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_379
timestamp 1556798218
transform 1 0 3704 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_378
timestamp 1556798218
transform -1 0 3800 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_377
timestamp 1556798218
transform 1 0 3800 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_427
timestamp 1556798218
transform 1 0 3848 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_130
timestamp 1556798218
transform -1 0 3944 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_383
timestamp 1556798218
transform 1 0 3944 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_384
timestamp 1556798218
transform -1 0 4072 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_131
timestamp 1556798218
transform -1 0 4136 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_163
timestamp 1556798218
transform 1 0 4136 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_425
timestamp 1556798218
transform -1 0 4216 0 -1 1010
box 0 0 32 200
use BUFX2  BUFX2_83
timestamp 1556798218
transform -1 0 4264 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_8
timestamp 1556798218
transform 1 0 4264 0 -1 1010
box 0 0 48 200
use XNOR2X1  XNOR2X1_62
timestamp 1556798218
transform 1 0 4312 0 -1 1010
box 0 0 112 200
use NAND2X1  NAND2X1_423
timestamp 1556798218
transform 1 0 4424 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_188
timestamp 1556798218
transform -1 0 4520 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_145
timestamp 1556798218
transform -1 0 4600 0 -1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_427
timestamp 1556798218
transform 1 0 4600 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_426
timestamp 1556798218
transform -1 0 4696 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_129
timestamp 1556798218
transform 1 0 4696 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_442
timestamp 1556798218
transform -1 0 4808 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_2_0
timestamp 1556798218
transform -1 0 4824 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1556798218
transform -1 0 4840 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_2
timestamp 1556798218
transform -1 0 4856 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_21
timestamp 1556798218
transform -1 0 4904 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_144
timestamp 1556798218
transform -1 0 4984 0 -1 1010
box 0 0 80 200
use INVX1  INVX1_489
timestamp 1556798218
transform 1 0 4984 0 -1 1010
box 0 0 32 200
use INVX1  INVX1_486
timestamp 1556798218
transform 1 0 5016 0 -1 1010
box 0 0 32 200
use INVX1  INVX1_491
timestamp 1556798218
transform 1 0 5048 0 -1 1010
box 0 0 32 200
use AND2X2  AND2X2_111
timestamp 1556798218
transform 1 0 5080 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_187
timestamp 1556798218
transform 1 0 5144 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_488
timestamp 1556798218
transform -1 0 5224 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_144
timestamp 1556798218
transform -1 0 5416 0 -1 1010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_142
timestamp 1556798218
transform 1 0 5416 0 -1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_199
timestamp 1556798218
transform 1 0 5608 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_224
timestamp 1556798218
transform -1 0 5720 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_242
timestamp 1556798218
transform -1 0 5752 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_147
timestamp 1556798218
transform 1 0 5752 0 -1 1010
box 0 0 192 200
use BUFX2  BUFX2_17
timestamp 1556798218
transform -1 0 5992 0 -1 1010
box 0 0 48 200
use CLKBUF1  CLKBUF1_31
timestamp 1556798218
transform -1 0 6136 0 -1 1010
box 0 0 144 200
use OAI21X1  OAI21X1_212
timestamp 1556798218
transform -1 0 6200 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_216
timestamp 1556798218
transform 1 0 6200 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_217
timestamp 1556798218
transform 1 0 6248 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_16
timestamp 1556798218
transform 1 0 6296 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_3_0
timestamp 1556798218
transform 1 0 6344 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_1
timestamp 1556798218
transform 1 0 6360 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_2
timestamp 1556798218
transform 1 0 6376 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_222
timestamp 1556798218
transform 1 0 6392 0 -1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_85
timestamp 1556798218
transform -1 0 6472 0 -1 1010
box 0 0 48 200
use XNOR2X1  XNOR2X1_28
timestamp 1556798218
transform -1 0 6584 0 -1 1010
box 0 0 112 200
use AOI21X1  AOI21X1_33
timestamp 1556798218
transform 1 0 6584 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_210
timestamp 1556798218
transform -1 0 6712 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_140
timestamp 1556798218
transform 1 0 6712 0 -1 1010
box 0 0 192 200
use INVX1  INVX1_226
timestamp 1556798218
transform -1 0 6936 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_181
timestamp 1556798218
transform 1 0 6936 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_57
timestamp 1556798218
transform 1 0 6984 0 -1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_73
timestamp 1556798218
transform -1 0 7112 0 -1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_117
timestamp 1556798218
transform -1 0 7304 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_171
timestamp 1556798218
transform -1 0 7368 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_60
timestamp 1556798218
transform -1 0 7432 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_179
timestamp 1556798218
transform 1 0 7432 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_61
timestamp 1556798218
transform -1 0 7544 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_173
timestamp 1556798218
transform -1 0 7608 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_267
timestamp 1556798218
transform -1 0 7800 0 -1 1010
box 0 0 192 200
use INVX1  INVX1_452
timestamp 1556798218
transform 1 0 7800 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_406
timestamp 1556798218
transform 1 0 7832 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_125
timestamp 1556798218
transform -1 0 8088 0 -1 1010
box 0 0 192 200
use AND2X2  AND2X2_8
timestamp 1556798218
transform 1 0 8088 0 -1 1010
box 0 0 64 200
use FILL  FILL_5_1
timestamp 1556798218
transform -1 0 8168 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_367
timestamp 1556798218
transform 1 0 8 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_368
timestamp 1556798218
transform -1 0 136 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_357
timestamp 1556798218
transform -1 0 184 0 1 610
box 0 0 48 200
use INVX1  INVX1_405
timestamp 1556798218
transform -1 0 216 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_359
timestamp 1556798218
transform 1 0 216 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_124
timestamp 1556798218
transform -1 0 328 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_120
timestamp 1556798218
transform -1 0 408 0 1 610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_245
timestamp 1556798218
transform 1 0 408 0 1 610
box 0 0 192 200
use INVX1  INVX1_165
timestamp 1556798218
transform -1 0 632 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_103
timestamp 1556798218
transform 1 0 632 0 1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_218
timestamp 1556798218
transform 1 0 824 0 1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_219
timestamp 1556798218
transform 1 0 1016 0 1 610
box 0 0 192 200
use INVX1  INVX1_368
timestamp 1556798218
transform -1 0 1240 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_132
timestamp 1556798218
transform -1 0 1288 0 1 610
box 0 0 48 200
use INVX1  INVX1_103
timestamp 1556798218
transform 1 0 1288 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_48
timestamp 1556798218
transform -1 0 1368 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_39
timestamp 1556798218
transform 1 0 1368 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_40
timestamp 1556798218
transform 1 0 1432 0 1 610
box 0 0 64 200
use INVX1  INVX1_108
timestamp 1556798218
transform 1 0 1496 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_105
timestamp 1556798218
transform 1 0 1528 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_49
timestamp 1556798218
transform 1 0 1592 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_35
timestamp 1556798218
transform -1 0 1720 0 1 610
box 0 0 80 200
use FILL  FILL_3_0_0
timestamp 1556798218
transform -1 0 1736 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1556798218
transform -1 0 1752 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_2
timestamp 1556798218
transform -1 0 1768 0 1 610
box 0 0 16 200
use OAI21X1  OAI21X1_107
timestamp 1556798218
transform -1 0 1832 0 1 610
box 0 0 64 200
use INVX1  INVX1_109
timestamp 1556798218
transform -1 0 1864 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_71
timestamp 1556798218
transform 1 0 1864 0 1 610
box 0 0 192 200
use CLKBUF1  CLKBUF1_15
timestamp 1556798218
transform 1 0 2056 0 1 610
box 0 0 144 200
use INVX1  INVX1_140
timestamp 1556798218
transform 1 0 2200 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_132
timestamp 1556798218
transform 1 0 2232 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_133
timestamp 1556798218
transform -1 0 2360 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_49
timestamp 1556798218
transform -1 0 2424 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_136
timestamp 1556798218
transform 1 0 2424 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_144
timestamp 1556798218
transform 1 0 2488 0 1 610
box 0 0 48 200
use INVX1  INVX1_139
timestamp 1556798218
transform -1 0 2568 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_60
timestamp 1556798218
transform 1 0 2568 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_44
timestamp 1556798218
transform -1 0 2696 0 1 610
box 0 0 80 200
use AOI22X1  AOI22X1_45
timestamp 1556798218
transform 1 0 2696 0 1 610
box 0 0 80 200
use OAI21X1  OAI21X1_134
timestamp 1556798218
transform 1 0 2776 0 1 610
box 0 0 64 200
use INVX1  INVX1_143
timestamp 1556798218
transform 1 0 2840 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_135
timestamp 1556798218
transform 1 0 2872 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_90
timestamp 1556798218
transform -1 0 3128 0 1 610
box 0 0 192 200
use CLKBUF1  CLKBUF1_33
timestamp 1556798218
transform 1 0 3128 0 1 610
box 0 0 144 200
use FILL  FILL_3_1_0
timestamp 1556798218
transform -1 0 3288 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1556798218
transform -1 0 3304 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_2
timestamp 1556798218
transform -1 0 3320 0 1 610
box 0 0 16 200
use NAND3X1  NAND3X1_109
timestamp 1556798218
transform -1 0 3384 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_129
timestamp 1556798218
transform 1 0 3384 0 1 610
box 0 0 48 200
use INVX1  INVX1_348
timestamp 1556798218
transform -1 0 3464 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_213
timestamp 1556798218
transform 1 0 3464 0 1 610
box 0 0 192 200
use BUFX2  BUFX2_115
timestamp 1556798218
transform -1 0 3704 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_375
timestamp 1556798218
transform -1 0 3752 0 1 610
box 0 0 48 200
use AND2X2  AND2X2_102
timestamp 1556798218
transform -1 0 3816 0 1 610
box 0 0 64 200
use INVX1  INVX1_429
timestamp 1556798218
transform 1 0 3816 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_385
timestamp 1556798218
transform -1 0 3912 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_62
timestamp 1556798218
transform 1 0 3912 0 1 610
box 0 0 64 200
use XNOR2X1  XNOR2X1_57
timestamp 1556798218
transform -1 0 4088 0 1 610
box 0 0 112 200
use OAI21X1  OAI21X1_387
timestamp 1556798218
transform 1 0 4088 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_376
timestamp 1556798218
transform -1 0 4200 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_116
timestamp 1556798218
transform -1 0 4248 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_4
timestamp 1556798218
transform 1 0 4248 0 1 610
box 0 0 48 200
use AND2X2  AND2X2_51
timestamp 1556798218
transform 1 0 4296 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_257
timestamp 1556798218
transform 1 0 4360 0 1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_109
timestamp 1556798218
transform -1 0 4744 0 1 610
box 0 0 192 200
use FILL  FILL_3_2_0
timestamp 1556798218
transform 1 0 4744 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1556798218
transform 1 0 4760 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_2
timestamp 1556798218
transform 1 0 4776 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_291
timestamp 1556798218
transform 1 0 4792 0 1 610
box 0 0 192 200
use INVX1  INVX1_494
timestamp 1556798218
transform -1 0 5016 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_434
timestamp 1556798218
transform 1 0 5016 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_433
timestamp 1556798218
transform 1 0 5080 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_143
timestamp 1556798218
transform -1 0 5224 0 1 610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_286
timestamp 1556798218
transform -1 0 5416 0 1 610
box 0 0 192 200
use AND2X2  AND2X2_11
timestamp 1556798218
transform 1 0 5416 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_223
timestamp 1556798218
transform 1 0 5480 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_436
timestamp 1556798218
transform -1 0 5592 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_149
timestamp 1556798218
transform 1 0 5592 0 1 610
box 0 0 192 200
use AND2X2  AND2X2_62
timestamp 1556798218
transform 1 0 5784 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_73
timestamp 1556798218
transform -1 0 5928 0 1 610
box 0 0 80 200
use NAND2X1  NAND2X1_227
timestamp 1556798218
transform 1 0 5928 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_226
timestamp 1556798218
transform -1 0 6024 0 1 610
box 0 0 48 200
use INVX1  INVX1_487
timestamp 1556798218
transform -1 0 6056 0 1 610
box 0 0 32 200
use INVX1  INVX1_206
timestamp 1556798218
transform 1 0 6056 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_287
timestamp 1556798218
transform 1 0 6088 0 1 610
box 0 0 192 200
use AND2X2  AND2X2_56
timestamp 1556798218
transform -1 0 6344 0 1 610
box 0 0 64 200
use FILL  FILL_3_3_0
timestamp 1556798218
transform 1 0 6344 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_1
timestamp 1556798218
transform 1 0 6360 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_2
timestamp 1556798218
transform 1 0 6376 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_194
timestamp 1556798218
transform 1 0 6392 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_196
timestamp 1556798218
transform 1 0 6440 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_198
timestamp 1556798218
transform 1 0 6488 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_197
timestamp 1556798218
transform -1 0 6584 0 1 610
box 0 0 48 200
use INVX1  INVX1_203
timestamp 1556798218
transform 1 0 6584 0 1 610
box 0 0 32 200
use XNOR2X1  XNOR2X1_25
timestamp 1556798218
transform -1 0 6728 0 1 610
box 0 0 112 200
use INVX1  INVX1_205
timestamp 1556798218
transform -1 0 6760 0 1 610
box 0 0 32 200
use AOI21X1  AOI21X1_30
timestamp 1556798218
transform 1 0 6760 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_128
timestamp 1556798218
transform 1 0 6824 0 1 610
box 0 0 192 200
use AND2X2  AND2X2_53
timestamp 1556798218
transform -1 0 7080 0 1 610
box 0 0 64 200
use BUFX2  BUFX2_107
timestamp 1556798218
transform -1 0 7128 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_110
timestamp 1556798218
transform -1 0 7176 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_166
timestamp 1556798218
transform -1 0 7224 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_67
timestamp 1556798218
transform -1 0 7272 0 1 610
box 0 0 48 200
use INVX1  INVX1_185
timestamp 1556798218
transform 1 0 7272 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_172
timestamp 1556798218
transform 1 0 7304 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_177
timestamp 1556798218
transform -1 0 7416 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_108
timestamp 1556798218
transform 1 0 7416 0 1 610
box 0 0 48 200
use INVX1  INVX1_184
timestamp 1556798218
transform -1 0 7496 0 1 610
box 0 0 32 200
use AOI21X1  AOI21X1_27
timestamp 1556798218
transform 1 0 7496 0 1 610
box 0 0 64 200
use XNOR2X1  XNOR2X1_22
timestamp 1556798218
transform -1 0 7672 0 1 610
box 0 0 112 200
use INVX1  INVX1_194
timestamp 1556798218
transform 1 0 7672 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_76
timestamp 1556798218
transform -1 0 7752 0 1 610
box 0 0 48 200
use INVX1  INVX1_284
timestamp 1556798218
transform -1 0 7784 0 1 610
box 0 0 32 200
use BUFX2  BUFX2_109
timestamp 1556798218
transform 1 0 7784 0 1 610
box 0 0 48 200
use INVX1  INVX1_195
timestamp 1556798218
transform 1 0 7832 0 1 610
box 0 0 32 200
use XNOR2X1  XNOR2X1_24
timestamp 1556798218
transform 1 0 7864 0 1 610
box 0 0 112 200
use NAND2X1  NAND2X1_190
timestamp 1556798218
transform -1 0 8024 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_65
timestamp 1556798218
transform 1 0 8024 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_183
timestamp 1556798218
transform 1 0 8088 0 1 610
box 0 0 64 200
use FILL  FILL_4_1
timestamp 1556798218
transform 1 0 8152 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_242
timestamp 1556798218
transform -1 0 200 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_361
timestamp 1556798218
transform 1 0 200 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_360
timestamp 1556798218
transform -1 0 296 0 -1 610
box 0 0 48 200
use INVX1  INVX1_407
timestamp 1556798218
transform -1 0 328 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_152
timestamp 1556798218
transform -1 0 376 0 -1 610
box 0 0 48 200
use AOI22X1  AOI22X1_121
timestamp 1556798218
transform -1 0 456 0 -1 610
box 0 0 80 200
use INVX1  INVX1_145
timestamp 1556798218
transform -1 0 488 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_370
timestamp 1556798218
transform -1 0 552 0 -1 610
box 0 0 64 200
use INVX1  INVX1_410
timestamp 1556798218
transform -1 0 584 0 -1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_243
timestamp 1556798218
transform 1 0 584 0 -1 610
box 0 0 192 200
use CLKBUF1  CLKBUF1_27
timestamp 1556798218
transform -1 0 920 0 -1 610
box 0 0 144 200
use CLKBUF1  CLKBUF1_43
timestamp 1556798218
transform 1 0 920 0 -1 610
box 0 0 144 200
use DFFPOSX1  DFFPOSX1_73
timestamp 1556798218
transform 1 0 1064 0 -1 610
box 0 0 192 200
use INVX1  INVX1_152
timestamp 1556798218
transform 1 0 1256 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_63
timestamp 1556798218
transform -1 0 1336 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_70
timestamp 1556798218
transform 1 0 1336 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_148
timestamp 1556798218
transform 1 0 1528 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_138
timestamp 1556798218
transform 1 0 1576 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_149
timestamp 1556798218
transform 1 0 1640 0 -1 610
box 0 0 48 200
use FILL  FILL_2_0_0
timestamp 1556798218
transform -1 0 1704 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1556798218
transform -1 0 1720 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_2
timestamp 1556798218
transform -1 0 1736 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_99
timestamp 1556798218
transform -1 0 1928 0 -1 610
box 0 0 192 200
use INVX1  INVX1_158
timestamp 1556798218
transform 1 0 1928 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_150
timestamp 1556798218
transform 1 0 1960 0 -1 610
box 0 0 64 200
use BUFX2  BUFX2_49
timestamp 1556798218
transform 1 0 2024 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_46
timestamp 1556798218
transform 1 0 2072 0 -1 610
box 0 0 48 200
use XNOR2X1  XNOR2X1_16
timestamp 1556798218
transform -1 0 2232 0 -1 610
box 0 0 112 200
use INVX1  INVX1_141
timestamp 1556798218
transform 1 0 2232 0 -1 610
box 0 0 32 200
use AND2X2  AND2X2_46
timestamp 1556798218
transform 1 0 2264 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_48
timestamp 1556798218
transform 1 0 2328 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_21
timestamp 1556798218
transform 1 0 2392 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_92
timestamp 1556798218
transform 1 0 2456 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_145
timestamp 1556798218
transform 1 0 2648 0 -1 610
box 0 0 48 200
use INVX1  INVX1_441
timestamp 1556798218
transform -1 0 2728 0 -1 610
box 0 0 32 200
use INVX1  INVX1_142
timestamp 1556798218
transform -1 0 2760 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_167
timestamp 1556798218
transform 1 0 2760 0 -1 610
box 0 0 48 200
use INVX1  INVX1_439
timestamp 1556798218
transform 1 0 2808 0 -1 610
box 0 0 32 200
use NAND2X1  NAND2X1_143
timestamp 1556798218
transform 1 0 2840 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_118
timestamp 1556798218
transform -1 0 2936 0 -1 610
box 0 0 48 200
use CLKBUF1  CLKBUF1_10
timestamp 1556798218
transform -1 0 3080 0 -1 610
box 0 0 144 200
use BUFX2  BUFX2_121
timestamp 1556798218
transform 1 0 3080 0 -1 610
box 0 0 48 200
use INVX1  INVX1_369
timestamp 1556798218
transform 1 0 3128 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_135
timestamp 1556798218
transform -1 0 3208 0 -1 610
box 0 0 48 200
use FILL  FILL_2_1_0
timestamp 1556798218
transform 1 0 3208 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1556798218
transform 1 0 3224 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_2
timestamp 1556798218
transform 1 0 3240 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_225
timestamp 1556798218
transform 1 0 3256 0 -1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_254
timestamp 1556798218
transform 1 0 3448 0 -1 610
box 0 0 192 200
use INVX1  INVX1_430
timestamp 1556798218
transform 1 0 3640 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_386
timestamp 1556798218
transform 1 0 3672 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_256
timestamp 1556798218
transform -1 0 3928 0 -1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_107
timestamp 1556798218
transform -1 0 4120 0 -1 610
box 0 0 192 200
use INVX1  INVX1_172
timestamp 1556798218
transform 1 0 4120 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_162
timestamp 1556798218
transform 1 0 4152 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_7
timestamp 1556798218
transform 1 0 4216 0 -1 610
box 0 0 48 200
use INVX1  INVX1_171
timestamp 1556798218
transform 1 0 4264 0 -1 610
box 0 0 32 200
use NAND2X1  NAND2X1_167
timestamp 1556798218
transform 1 0 4296 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_160
timestamp 1556798218
transform 1 0 4344 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_106
timestamp 1556798218
transform -1 0 4600 0 -1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_289
timestamp 1556798218
transform 1 0 4600 0 -1 610
box 0 0 192 200
use BUFX2  BUFX2_134
timestamp 1556798218
transform 1 0 4792 0 -1 610
box 0 0 48 200
use FILL  FILL_2_2_0
timestamp 1556798218
transform 1 0 4840 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1556798218
transform 1 0 4856 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_2
timestamp 1556798218
transform 1 0 4872 0 -1 610
box 0 0 16 200
use INVX1  INVX1_482
timestamp 1556798218
transform 1 0 4888 0 -1 610
box 0 0 32 200
use INVX1  INVX1_483
timestamp 1556798218
transform 1 0 4920 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_186
timestamp 1556798218
transform 1 0 4952 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_418
timestamp 1556798218
transform 1 0 5000 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_420
timestamp 1556798218
transform 1 0 5048 0 -1 610
box 0 0 48 200
use AOI22X1  AOI22X1_142
timestamp 1556798218
transform -1 0 5176 0 -1 610
box 0 0 80 200
use NAND2X1  NAND2X1_421
timestamp 1556798218
transform 1 0 5176 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_422
timestamp 1556798218
transform -1 0 5272 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_146
timestamp 1556798218
transform 1 0 5272 0 -1 610
box 0 0 192 200
use INVX1  INVX1_241
timestamp 1556798218
transform 1 0 5464 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_222
timestamp 1556798218
transform 1 0 5496 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_221
timestamp 1556798218
transform -1 0 5624 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_225
timestamp 1556798218
transform 1 0 5624 0 -1 610
box 0 0 48 200
use AOI22X1  AOI22X1_72
timestamp 1556798218
transform -1 0 5752 0 -1 610
box 0 0 80 200
use INVX1  INVX1_239
timestamp 1556798218
transform -1 0 5784 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_90
timestamp 1556798218
transform -1 0 5832 0 -1 610
box 0 0 48 200
use INVX1  INVX1_238
timestamp 1556798218
transform -1 0 5864 0 -1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_126
timestamp 1556798218
transform 1 0 5864 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_191
timestamp 1556798218
transform 1 0 6056 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_190
timestamp 1556798218
transform -1 0 6184 0 -1 610
box 0 0 64 200
use INVX1  INVX1_202
timestamp 1556798218
transform 1 0 6184 0 -1 610
box 0 0 32 200
use AOI22X1  AOI22X1_63
timestamp 1556798218
transform -1 0 6296 0 -1 610
box 0 0 80 200
use NOR2X1  NOR2X1_79
timestamp 1556798218
transform 1 0 6296 0 -1 610
box 0 0 48 200
use FILL  FILL_2_3_0
timestamp 1556798218
transform 1 0 6344 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_1
timestamp 1556798218
transform 1 0 6360 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_2
timestamp 1556798218
transform 1 0 6376 0 -1 610
box 0 0 16 200
use AOI22X1  AOI22X1_62
timestamp 1556798218
transform 1 0 6392 0 -1 610
box 0 0 80 200
use NAND3X1  NAND3X1_66
timestamp 1556798218
transform -1 0 6536 0 -1 610
box 0 0 64 200
use INVX1  INVX1_204
timestamp 1556798218
transform -1 0 6568 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_188
timestamp 1556798218
transform 1 0 6568 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_189
timestamp 1556798218
transform -1 0 6696 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_67
timestamp 1556798218
transform -1 0 6760 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_195
timestamp 1556798218
transform 1 0 6760 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_192
timestamp 1556798218
transform 1 0 6808 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_78
timestamp 1556798218
transform 1 0 6872 0 -1 610
box 0 0 48 200
use INVX1  INVX1_201
timestamp 1556798218
transform -1 0 6952 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_63
timestamp 1556798218
transform -1 0 7016 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_177
timestamp 1556798218
transform 1 0 7016 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_185
timestamp 1556798218
transform -1 0 7128 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_180
timestamp 1556798218
transform 1 0 7128 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_74
timestamp 1556798218
transform 1 0 7192 0 -1 610
box 0 0 48 200
use INVX1  INVX1_187
timestamp 1556798218
transform -1 0 7272 0 -1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_114
timestamp 1556798218
transform -1 0 7464 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_165
timestamp 1556798218
transform -1 0 7512 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_116
timestamp 1556798218
transform -1 0 7704 0 -1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_124
timestamp 1556798218
transform 1 0 7704 0 -1 610
box 0 0 192 200
use INVX1  INVX1_198
timestamp 1556798218
transform 1 0 7896 0 -1 610
box 0 0 32 200
use AOI21X1  AOI21X1_29
timestamp 1556798218
transform 1 0 7928 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_186
timestamp 1556798218
transform -1 0 8056 0 -1 610
box 0 0 64 200
use INVX1  INVX1_197
timestamp 1556798218
transform 1 0 8056 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_182
timestamp 1556798218
transform -1 0 8152 0 -1 610
box 0 0 64 200
use FILL  FILL_3_1
timestamp 1556798218
transform -1 0 8168 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_97
timestamp 1556798218
transform -1 0 200 0 1 210
box 0 0 192 200
use NAND3X1  NAND3X1_51
timestamp 1556798218
transform -1 0 264 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_143
timestamp 1556798218
transform 1 0 264 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_50
timestamp 1556798218
transform 1 0 328 0 1 210
box 0 0 64 200
use INVX1  INVX1_148
timestamp 1556798218
transform 1 0 392 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_61
timestamp 1556798218
transform 1 0 424 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_153
timestamp 1556798218
transform 1 0 472 0 1 210
box 0 0 48 200
use AOI21X1  AOI21X1_22
timestamp 1556798218
transform -1 0 584 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_154
timestamp 1556798218
transform -1 0 632 0 1 210
box 0 0 48 200
use INVX1  INVX1_149
timestamp 1556798218
transform -1 0 664 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_96
timestamp 1556798218
transform 1 0 664 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_144
timestamp 1556798218
transform -1 0 920 0 1 210
box 0 0 64 200
use INVX1  INVX1_151
timestamp 1556798218
transform -1 0 952 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_95
timestamp 1556798218
transform 1 0 952 0 1 210
box 0 0 192 200
use BUFX2  BUFX2_47
timestamp 1556798218
transform -1 0 1192 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_54
timestamp 1556798218
transform 1 0 1192 0 1 210
box 0 0 48 200
use XNOR2X1  XNOR2X1_18
timestamp 1556798218
transform 1 0 1240 0 1 210
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_101
timestamp 1556798218
transform 1 0 1352 0 1 210
box 0 0 192 200
use NAND3X1  NAND3X1_53
timestamp 1556798218
transform 1 0 1544 0 1 210
box 0 0 64 200
use INVX1  INVX1_154
timestamp 1556798218
transform 1 0 1608 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_145
timestamp 1556798218
transform -1 0 1704 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_146
timestamp 1556798218
transform -1 0 1768 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1556798218
transform -1 0 1784 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1556798218
transform -1 0 1800 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_2
timestamp 1556798218
transform -1 0 1816 0 1 210
box 0 0 16 200
use AOI22X1  AOI22X1_48
timestamp 1556798218
transform -1 0 1896 0 1 210
box 0 0 80 200
use NAND2X1  NAND2X1_158
timestamp 1556798218
transform 1 0 1896 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_98
timestamp 1556798218
transform -1 0 2136 0 1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_263
timestamp 1556798218
transform 1 0 2136 0 1 210
box 0 0 192 200
use INVX1  INVX1_445
timestamp 1556798218
transform 1 0 2328 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_400
timestamp 1556798218
transform 1 0 2360 0 1 210
box 0 0 64 200
use INVX1  INVX1_442
timestamp 1556798218
transform 1 0 2424 0 1 210
box 0 0 32 200
use AOI22X1  AOI22X1_130
timestamp 1556798218
transform -1 0 2536 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_399
timestamp 1556798218
transform 1 0 2536 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_387
timestamp 1556798218
transform -1 0 2648 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_395
timestamp 1556798218
transform 1 0 2648 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_396
timestamp 1556798218
transform -1 0 2776 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_388
timestamp 1556798218
transform -1 0 2824 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_135
timestamp 1556798218
transform 1 0 2824 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_134
timestamp 1556798218
transform 1 0 2888 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_168
timestamp 1556798218
transform -1 0 3000 0 1 210
box 0 0 48 200
use AOI22X1  AOI22X1_131
timestamp 1556798218
transform -1 0 3080 0 1 210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_265
timestamp 1556798218
transform 1 0 3080 0 1 210
box 0 0 192 200
use FILL  FILL_1_1_0
timestamp 1556798218
transform 1 0 3272 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1556798218
transform 1 0 3288 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_2
timestamp 1556798218
transform 1 0 3304 0 1 210
box 0 0 16 200
use NAND3X1  NAND3X1_115
timestamp 1556798218
transform 1 0 3320 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_339
timestamp 1556798218
transform -1 0 3448 0 1 210
box 0 0 64 200
use INVX1  INVX1_371
timestamp 1556798218
transform 1 0 3448 0 1 210
box 0 0 32 200
use NAND2X1  NAND2X1_330
timestamp 1556798218
transform 1 0 3480 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_336
timestamp 1556798218
transform 1 0 3528 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_335
timestamp 1556798218
transform -1 0 3656 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_114
timestamp 1556798218
transform 1 0 3656 0 1 210
box 0 0 64 200
use INVX1  INVX1_370
timestamp 1556798218
transform -1 0 3752 0 1 210
box 0 0 32 200
use AND2X2  AND2X2_86
timestamp 1556798218
transform 1 0 3752 0 1 210
box 0 0 64 200
use INVX1  INVX1_374
timestamp 1556798218
transform 1 0 3816 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_338
timestamp 1556798218
transform 1 0 3848 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_337
timestamp 1556798218
transform 1 0 3912 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_111
timestamp 1556798218
transform -1 0 4056 0 1 210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_222
timestamp 1556798218
transform 1 0 4056 0 1 210
box 0 0 192 200
use BUFX2  BUFX2_85
timestamp 1556798218
transform 1 0 4248 0 1 210
box 0 0 48 200
use AOI22X1  AOI22X1_53
timestamp 1556798218
transform 1 0 4296 0 1 210
box 0 0 80 200
use NOR2X1  NOR2X1_69
timestamp 1556798218
transform 1 0 4376 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_159
timestamp 1556798218
transform -1 0 4488 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_52
timestamp 1556798218
transform -1 0 4568 0 1 210
box 0 0 80 200
use INVX1  INVX1_170
timestamp 1556798218
transform 1 0 4568 0 1 210
box 0 0 32 200
use NAND3X1  NAND3X1_56
timestamp 1556798218
transform -1 0 4664 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_57
timestamp 1556798218
transform -1 0 4728 0 1 210
box 0 0 64 200
use XNOR2X1  XNOR2X1_20
timestamp 1556798218
transform -1 0 4840 0 1 210
box 0 0 112 200
use FILL  FILL_1_2_0
timestamp 1556798218
transform 1 0 4840 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1556798218
transform 1 0 4856 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_2
timestamp 1556798218
transform 1 0 4872 0 1 210
box 0 0 16 200
use INVX1  INVX1_166
timestamp 1556798218
transform 1 0 4888 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_68
timestamp 1556798218
transform -1 0 4968 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_431
timestamp 1556798218
transform 1 0 4968 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_432
timestamp 1556798218
transform -1 0 5096 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_147
timestamp 1556798218
transform -1 0 5160 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_419
timestamp 1556798218
transform -1 0 5208 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_146
timestamp 1556798218
transform 1 0 5208 0 1 210
box 0 0 64 200
use INVX1  INVX1_484
timestamp 1556798218
transform -1 0 5304 0 1 210
box 0 0 32 200
use XNOR2X1  XNOR2X1_65
timestamp 1556798218
transform -1 0 5416 0 1 210
box 0 0 112 200
use AND2X2  AND2X2_10
timestamp 1556798218
transform -1 0 5480 0 1 210
box 0 0 64 200
use INVX1  INVX1_236
timestamp 1556798218
transform 1 0 5480 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_89
timestamp 1556798218
transform -1 0 5560 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_76
timestamp 1556798218
transform -1 0 5624 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_77
timestamp 1556798218
transform 1 0 5624 0 1 210
box 0 0 64 200
use INVX1  INVX1_237
timestamp 1556798218
transform -1 0 5720 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_220
timestamp 1556798218
transform 1 0 5720 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_219
timestamp 1556798218
transform 1 0 5784 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_223
timestamp 1556798218
transform -1 0 5912 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_224
timestamp 1556798218
transform -1 0 5960 0 1 210
box 0 0 48 200
use CLKBUF1  CLKBUF1_4
timestamp 1556798218
transform -1 0 6104 0 1 210
box 0 0 144 200
use CLKBUF1  CLKBUF1_16
timestamp 1556798218
transform 1 0 6104 0 1 210
box 0 0 144 200
use OAI21X1  OAI21X1_193
timestamp 1556798218
transform -1 0 6312 0 1 210
box 0 0 64 200
use INVX1  INVX1_207
timestamp 1556798218
transform -1 0 6344 0 1 210
box 0 0 32 200
use FILL  FILL_1_3_0
timestamp 1556798218
transform -1 0 6360 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_1
timestamp 1556798218
transform -1 0 6376 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_2
timestamp 1556798218
transform -1 0 6392 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_129
timestamp 1556798218
transform -1 0 6584 0 1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_121
timestamp 1556798218
transform -1 0 6776 0 1 210
box 0 0 192 200
use INVX1  INVX1_188
timestamp 1556798218
transform -1 0 6808 0 1 210
box 0 0 32 200
use NAND2X1  NAND2X1_188
timestamp 1556798218
transform 1 0 6808 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_187
timestamp 1556798218
transform 1 0 6856 0 1 210
box 0 0 48 200
use INVX1  INVX1_190
timestamp 1556798218
transform -1 0 6936 0 1 210
box 0 0 32 200
use NAND3X1  NAND3X1_62
timestamp 1556798218
transform -1 0 7000 0 1 210
box 0 0 64 200
use INVX1  INVX1_189
timestamp 1556798218
transform 1 0 7000 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_176
timestamp 1556798218
transform 1 0 7032 0 1 210
box 0 0 64 200
use XNOR2X1  XNOR2X1_23
timestamp 1556798218
transform -1 0 7208 0 1 210
box 0 0 112 200
use AOI21X1  AOI21X1_28
timestamp 1556798218
transform 1 0 7208 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_120
timestamp 1556798218
transform 1 0 7272 0 1 210
box 0 0 192 200
use CLKBUF1  CLKBUF1_49
timestamp 1556798218
transform 1 0 7464 0 1 210
box 0 0 144 200
use INVX1  INVX1_199
timestamp 1556798218
transform -1 0 7640 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_185
timestamp 1556798218
transform 1 0 7640 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_189
timestamp 1556798218
transform -1 0 7752 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_184
timestamp 1556798218
transform -1 0 7816 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_191
timestamp 1556798218
transform 1 0 7816 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_192
timestamp 1556798218
transform -1 0 7912 0 1 210
box 0 0 48 200
use AOI22X1  AOI22X1_60
timestamp 1556798218
transform 1 0 7912 0 1 210
box 0 0 80 200
use AND2X2  AND2X2_55
timestamp 1556798218
transform 1 0 7992 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_77
timestamp 1556798218
transform -1 0 8104 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_137
timestamp 1556798218
transform 1 0 8104 0 1 210
box 0 0 48 200
use FILL  FILL_2_1
timestamp 1556798218
transform 1 0 8152 0 1 210
box 0 0 16 200
use AND2X2  AND2X2_5
timestamp 1556798218
transform 1 0 8 0 -1 210
box 0 0 64 200
use INVX1  INVX1_147
timestamp 1556798218
transform 1 0 72 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_139
timestamp 1556798218
transform -1 0 168 0 -1 210
box 0 0 64 200
use INVX1  INVX1_146
timestamp 1556798218
transform 1 0 168 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_140
timestamp 1556798218
transform -1 0 264 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_151
timestamp 1556798218
transform 1 0 264 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_152
timestamp 1556798218
transform 1 0 312 0 -1 210
box 0 0 48 200
use AOI22X1  AOI22X1_46
timestamp 1556798218
transform -1 0 440 0 -1 210
box 0 0 80 200
use NOR2X1  NOR2X1_62
timestamp 1556798218
transform -1 0 488 0 -1 210
box 0 0 48 200
use XNOR2X1  XNOR2X1_17
timestamp 1556798218
transform 1 0 488 0 -1 210
box 0 0 112 200
use AND2X2  AND2X2_47
timestamp 1556798218
transform 1 0 600 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_47
timestamp 1556798218
transform 1 0 664 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_141
timestamp 1556798218
transform 1 0 744 0 -1 210
box 0 0 64 200
use INVX1  INVX1_150
timestamp 1556798218
transform 1 0 808 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_150
timestamp 1556798218
transform 1 0 840 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_142
timestamp 1556798218
transform 1 0 888 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_94
timestamp 1556798218
transform -1 0 1144 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_131
timestamp 1556798218
transform -1 0 1192 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_100
timestamp 1556798218
transform -1 0 1384 0 -1 210
box 0 0 192 200
use AOI21X1  AOI21X1_23
timestamp 1556798218
transform 1 0 1384 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_149
timestamp 1556798218
transform -1 0 1512 0 -1 210
box 0 0 64 200
use INVX1  INVX1_156
timestamp 1556798218
transform 1 0 1512 0 -1 210
box 0 0 32 200
use NAND3X1  NAND3X1_52
timestamp 1556798218
transform -1 0 1608 0 -1 210
box 0 0 64 200
use INVX1  INVX1_153
timestamp 1556798218
transform 1 0 1608 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_156
timestamp 1556798218
transform -1 0 1688 0 -1 210
box 0 0 48 200
use INVX1  INVX1_155
timestamp 1556798218
transform -1 0 1720 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_157
timestamp 1556798218
transform 1 0 1720 0 -1 210
box 0 0 48 200
use FILL  FILL_0_0_0
timestamp 1556798218
transform -1 0 1784 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1556798218
transform -1 0 1800 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_2
timestamp 1556798218
transform -1 0 1816 0 -1 210
box 0 0 16 200
use NOR2X1  NOR2X1_64
timestamp 1556798218
transform -1 0 1864 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_147
timestamp 1556798218
transform 1 0 1864 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_159
timestamp 1556798218
transform -1 0 1976 0 -1 210
box 0 0 48 200
use AOI22X1  AOI22X1_49
timestamp 1556798218
transform -1 0 2056 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_148
timestamp 1556798218
transform -1 0 2120 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_155
timestamp 1556798218
transform -1 0 2168 0 -1 210
box 0 0 48 200
use INVX1  INVX1_157
timestamp 1556798218
transform -1 0 2200 0 -1 210
box 0 0 32 200
use AND2X2  AND2X2_48
timestamp 1556798218
transform -1 0 2264 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_7
timestamp 1556798218
transform -1 0 2328 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_264
timestamp 1556798218
transform -1 0 2520 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_386
timestamp 1556798218
transform 1 0 2520 0 -1 210
box 0 0 48 200
use AOI21X1  AOI21X1_64
timestamp 1556798218
transform -1 0 2632 0 -1 210
box 0 0 64 200
use XNOR2X1  XNOR2X1_59
timestamp 1556798218
transform -1 0 2744 0 -1 210
box 0 0 112 200
use INVX1  INVX1_440
timestamp 1556798218
transform -1 0 2776 0 -1 210
box 0 0 32 200
use INVX1  INVX1_443
timestamp 1556798218
transform 1 0 2776 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_389
timestamp 1556798218
transform -1 0 2856 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_385
timestamp 1556798218
transform -1 0 2904 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_397
timestamp 1556798218
transform 1 0 2904 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_398
timestamp 1556798218
transform -1 0 3032 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_262
timestamp 1556798218
transform -1 0 3224 0 -1 210
box 0 0 192 200
use INVX1  INVX1_444
timestamp 1556798218
transform -1 0 3256 0 -1 210
box 0 0 32 200
use FILL  FILL_0_1_0
timestamp 1556798218
transform -1 0 3272 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1556798218
transform -1 0 3288 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_2
timestamp 1556798218
transform -1 0 3304 0 -1 210
box 0 0 16 200
use XNOR2X1  XNOR2X1_49
timestamp 1556798218
transform -1 0 3416 0 -1 210
box 0 0 112 200
use AOI21X1  AOI21X1_54
timestamp 1556798218
transform -1 0 3480 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_224
timestamp 1556798218
transform 1 0 3480 0 -1 210
box 0 0 192 200
use INVX1  INVX1_373
timestamp 1556798218
transform -1 0 3704 0 -1 210
box 0 0 32 200
use INVX1  INVX1_372
timestamp 1556798218
transform -1 0 3736 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_331
timestamp 1556798218
transform 1 0 3736 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_329
timestamp 1556798218
transform 1 0 3784 0 -1 210
box 0 0 48 200
use AOI22X1  AOI22X1_110
timestamp 1556798218
transform -1 0 3912 0 -1 210
box 0 0 80 200
use NOR2X1  NOR2X1_136
timestamp 1556798218
transform -1 0 3960 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_332
timestamp 1556798218
transform 1 0 3960 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_333
timestamp 1556798218
transform -1 0 4056 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_340
timestamp 1556798218
transform -1 0 4120 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_223
timestamp 1556798218
transform 1 0 4120 0 -1 210
box 0 0 192 200
use INVX1  INVX1_375
timestamp 1556798218
transform -1 0 4344 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_171
timestamp 1556798218
transform 1 0 4344 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_170
timestamp 1556798218
transform -1 0 4440 0 -1 210
box 0 0 48 200
use INVX1  INVX1_169
timestamp 1556798218
transform -1 0 4472 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_169
timestamp 1556798218
transform -1 0 4520 0 -1 210
box 0 0 48 200
use INVX1  INVX1_167
timestamp 1556798218
transform -1 0 4552 0 -1 210
box 0 0 32 200
use INVX1  INVX1_168
timestamp 1556798218
transform 1 0 4552 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_157
timestamp 1556798218
transform 1 0 4584 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_158
timestamp 1556798218
transform -1 0 4712 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_168
timestamp 1556798218
transform -1 0 4760 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_161
timestamp 1556798218
transform 1 0 4760 0 -1 210
box 0 0 64 200
use FILL  FILL_0_2_0
timestamp 1556798218
transform 1 0 4824 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1556798218
transform 1 0 4840 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_2
timestamp 1556798218
transform 1 0 4856 0 -1 210
box 0 0 16 200
use AOI21X1  AOI21X1_25
timestamp 1556798218
transform 1 0 4872 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_108
timestamp 1556798218
transform -1 0 5128 0 -1 210
box 0 0 192 200
use INVX1  INVX1_485
timestamp 1556798218
transform 1 0 5128 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_435
timestamp 1556798218
transform 1 0 5160 0 -1 210
box 0 0 64 200
use INVX1  INVX1_481
timestamp 1556798218
transform 1 0 5224 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_185
timestamp 1556798218
transform -1 0 5304 0 -1 210
box 0 0 48 200
use AOI21X1  AOI21X1_70
timestamp 1556798218
transform -1 0 5368 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_288
timestamp 1556798218
transform -1 0 5560 0 -1 210
box 0 0 192 200
use INVX1  INVX1_240
timestamp 1556798218
transform 1 0 5560 0 -1 210
box 0 0 32 200
use XNOR2X1  XNOR2X1_30
timestamp 1556798218
transform -1 0 5704 0 -1 210
box 0 0 112 200
use AOI21X1  AOI21X1_35
timestamp 1556798218
transform 1 0 5704 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_148
timestamp 1556798218
transform -1 0 5960 0 -1 210
box 0 0 192 200
use AND2X2  AND2X2_3
timestamp 1556798218
transform 1 0 5960 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_127
timestamp 1556798218
transform 1 0 6024 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_118
timestamp 1556798218
transform 1 0 6216 0 -1 210
box 0 0 192 200
use FILL  FILL_0_3_0
timestamp 1556798218
transform 1 0 6408 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_1
timestamp 1556798218
transform 1 0 6424 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_2
timestamp 1556798218
transform 1 0 6440 0 -1 210
box 0 0 16 200
use AND2X2  AND2X2_54
timestamp 1556798218
transform 1 0 6456 0 -1 210
box 0 0 64 200
use INVX1  INVX1_192
timestamp 1556798218
transform 1 0 6520 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_179
timestamp 1556798218
transform 1 0 6552 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_184
timestamp 1556798218
transform 1 0 6616 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_178
timestamp 1556798218
transform -1 0 6728 0 -1 210
box 0 0 64 200
use INVX1  INVX1_191
timestamp 1556798218
transform 1 0 6728 0 -1 210
box 0 0 32 200
use AOI22X1  AOI22X1_59
timestamp 1556798218
transform -1 0 6840 0 -1 210
box 0 0 80 200
use NOR2X1  NOR2X1_75
timestamp 1556798218
transform 1 0 6840 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_186
timestamp 1556798218
transform 1 0 6888 0 -1 210
box 0 0 48 200
use AOI22X1  AOI22X1_58
timestamp 1556798218
transform -1 0 7016 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_181
timestamp 1556798218
transform -1 0 7080 0 -1 210
box 0 0 64 200
use INVX1  INVX1_193
timestamp 1556798218
transform -1 0 7112 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_119
timestamp 1556798218
transform -1 0 7304 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_182
timestamp 1556798218
transform 1 0 7304 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_183
timestamp 1556798218
transform 1 0 7352 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_175
timestamp 1556798218
transform 1 0 7400 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_123
timestamp 1556798218
transform -1 0 7656 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_122
timestamp 1556798218
transform 1 0 7656 0 -1 210
box 0 0 192 200
use INVX1  INVX1_200
timestamp 1556798218
transform 1 0 7848 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_193
timestamp 1556798218
transform 1 0 7880 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_187
timestamp 1556798218
transform 1 0 7928 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_61
timestamp 1556798218
transform -1 0 8072 0 -1 210
box 0 0 80 200
use NAND3X1  NAND3X1_64
timestamp 1556798218
transform 1 0 8072 0 -1 210
box 0 0 64 200
use FILL  FILL_1_1
timestamp 1556798218
transform -1 0 8152 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1556798218
transform -1 0 8168 0 -1 210
box 0 0 16 200
<< labels >>
flabel metal4 s 1736 0 1784 24 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 3272 0 3320 24 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 6205 5837 6211 5843 3 FreeSans 24 90 0 0 CLK
port 2 nsew
flabel metal2 s 2429 5837 2435 5843 3 FreeSans 24 90 0 0 RST_N
port 3 nsew
flabel metal2 s 4029 5837 4035 5843 3 FreeSans 24 90 0 0 request_put[0]
port 4 nsew
flabel metal2 s 2509 5837 2515 5843 3 FreeSans 24 90 0 0 request_put[1]
port 5 nsew
flabel metal2 s 2621 5837 2627 5843 3 FreeSans 24 90 0 0 request_put[2]
port 6 nsew
flabel metal2 s 2813 5837 2819 5843 3 FreeSans 24 90 0 0 request_put[3]
port 7 nsew
flabel metal2 s 3069 5837 3075 5843 3 FreeSans 24 90 0 0 request_put[4]
port 8 nsew
flabel metal2 s 3805 5837 3811 5843 3 FreeSans 24 90 0 0 request_put[5]
port 9 nsew
flabel metal2 s 3613 5837 3619 5843 3 FreeSans 24 90 0 0 request_put[6]
port 10 nsew
flabel metal2 s 4381 5837 4387 5843 3 FreeSans 24 90 0 0 EN_request_put
port 11 nsew
flabel metal3 s 8189 2497 8195 2503 3 FreeSans 24 0 0 0 EN_response_get
port 12 nsew
flabel metal2 s 3917 5837 3923 5843 3 FreeSans 24 90 0 0 RDY_request_put
port 13 nsew
flabel metal3 s 8189 297 8195 303 3 FreeSans 24 0 0 0 response_get[0]
port 14 nsew
flabel metal3 s 8189 3297 8195 3303 3 FreeSans 24 0 0 0 response_get[1]
port 15 nsew
flabel metal3 s 8189 1937 8195 1943 3 FreeSans 24 0 0 0 response_get[2]
port 16 nsew
flabel metal3 s 8189 3337 8195 3343 3 FreeSans 24 0 0 0 response_get[3]
port 17 nsew
flabel metal3 s 8189 1897 8195 1903 3 FreeSans 24 0 0 0 response_get[4]
port 18 nsew
flabel metal3 s 8189 2097 8195 2103 3 FreeSans 24 0 0 0 response_get[5]
port 19 nsew
flabel metal3 s 8189 2897 8195 2903 3 FreeSans 24 0 0 0 response_get[6]
port 20 nsew
flabel metal3 s 8189 5097 8195 5103 3 FreeSans 24 0 0 0 RDY_response_get
port 21 nsew
<< end >>
