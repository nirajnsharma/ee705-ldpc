* NGSPICE file created from mkLdpcCore.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

.subckt mkLdpcCore vdd gnd CLK RST_N request_put[0] request_put[1] request_put[2]
+ request_put[3] request_put[4] request_put[5] request_put[6] EN_request_put EN_response_get
+ RDY_request_put response_get[0] response_get[1] response_get[2] response_get[3]
+ response_get[4] response_get[5] response_get[6] RDY_response_get
XNAND2X1_376 BUFX2_116/Y INVX1_426/Y gnd OAI21X1_387/B vdd NAND2X1
XINVX1_624 INVX1_624/A gnd INVX1_624/Y vdd INVX1
XNOR2X1_62 AND2X2_5/B NOR2X1_62/B gnd NOR2X1_62/Y vdd NOR2X1
XOAI21X1_226 BUFX2_14/Y INVX1_244/Y OAI21X1_226/C gnd NAND3X1_79/C vdd OAI21X1
XNAND2X1_340 INVX1_378/A BUFX2_37/Y gnd NAND2X1_340/Y vdd NAND2X1
XCLKBUF1_50 BUFX2_3/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XINVX1_588 INVX1_588/A gnd INVX1_588/Y vdd INVX1
XNAND3X1_172 BUFX2_124/Y INVX1_575/Y INVX1_576/Y gnd NAND3X1_172/Y vdd NAND3X1
XOAI21X1_190 INVX1_202/Y INVX1_205/Y AOI22X1_63/C gnd OAI21X1_191/C vdd OAI21X1
XNOR2X1_26 AOI22X1_9/C INVX1_39/A gnd NOR2X1_26/Y vdd NOR2X1
XFILL_12_2_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_223 gnd INVX1_572/Y gnd NOR2X1_223/Y vdd NOR2X1
XNAND2X1_304 BUFX2_26/Y INVX1_338/A gnd OAI21X1_308/B vdd NAND2X1
XNAND3X1_136 BUFX2_113/Y INVX1_449/Y INVX1_450/Y gnd NAND3X1_136/Y vdd NAND3X1
XINVX1_552 BUFX2_97/Y gnd INVX1_552/Y vdd INVX1
XCLKBUF1_14 BUFX2_3/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XBUFX2_137 BUFX2_137/A gnd response_get[0] vdd BUFX2
XNOR2X1_187 gnd INVX1_488/Y gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_154 INVX1_164/Y NAND2X1_160/Y OAI21X1_153/Y gnd OAI21X1_154/Y vdd OAI21X1
XNAND2X1_268 INVX1_308/A INVX1_331/A gnd NOR2X1_106/B vdd NAND2X1
XFILL_0_0_2 gnd vdd FILL
XBUFX2_101 BUFX2_98/A gnd INVX1_475/A vdd BUFX2
XDFFPOSX1_334 AOI22X1_167/C CLKBUF1_23/Y OAI21X1_506/Y gnd vdd DFFPOSX1
XNAND3X1_100 INVX1_582/A INVX1_323/Y INVX1_324/Y gnd NAND3X1_100/Y vdd NAND3X1
XINVX1_516 BUFX2_33/Y gnd INVX1_516/Y vdd INVX1
XOAI21X1_118 INVX1_119/Y OAI21X1_118/B NOR2X1_52/Y gnd AOI21X1_18/C vdd OAI21X1
XXNOR2X1_61 AND2X2_9/Y BUFX2_112/Y gnd XNOR2X1_61/Y vdd XNOR2X1
XNOR2X1_151 gnd INVX1_404/Y gnd NOR2X1_151/Y vdd NOR2X1
XNAND2X1_232 INVX1_247/A NAND2X1_231/Y gnd AOI22X1_75/A vdd NAND2X1
XDFFPOSX1_298 AOI22X1_149/C CLKBUF1_12/Y OAI21X1_452/Y gnd vdd DFFPOSX1
XINVX1_480 INVX1_480/A gnd INVX1_480/Y vdd INVX1
XXNOR2X1_25 INVX1_204/A INVX1_484/A gnd XNOR2X1_25/Y vdd XNOR2X1
XNOR2X1_115 gnd INVX1_320/Y gnd NOR2X1_115/Y vdd NOR2X1
XNAND2X1_196 INVX1_484/A INVX1_205/Y gnd AOI22X1_62/D vdd NAND2X1
XINVX1_444 INVX1_444/A gnd INVX1_444/Y vdd INVX1
XDFFPOSX1_262 OAI21X1_397/C CLKBUF1_10/Y OAI21X1_398/Y gnd vdd DFFPOSX1
XFILL_21_0_0 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XBUFX2_97 BUFX2_96/A gnd BUFX2_97/Y vdd BUFX2
XFILL_19_2_1 gnd vdd FILL
XNAND2X1_160 INVX1_160/A INVX1_163/A gnd NAND2X1_160/Y vdd NAND2X1
XDFFPOSX1_226 AOI22X1_113/C CLKBUF1_41/Y OAI21X1_344/Y gnd vdd DFFPOSX1
XINVX1_408 AND2X2_5/A gnd INVX1_408/Y vdd INVX1
XAOI21X1_58 INVX1_401/Y AOI21X1_58/B AOI21X1_58/C gnd AOI21X1_58/Y vdd AOI21X1
XBUFX2_61 BUFX2_65/A gnd BUFX2_61/Y vdd BUFX2
XNAND2X1_124 AND2X2_4/B INVX1_106/A gnd NAND2X1_124/Y vdd NAND2X1
XFILL_7_0_2 gnd vdd FILL
XAOI21X1_22 INVX1_149/Y XNOR2X1_17/Y AOI21X1_22/C gnd AOI21X1_22/Y vdd AOI21X1
XFILL_9_1 gnd vdd FILL
XDFFPOSX1_190 AOI22X1_95/C CLKBUF1_32/Y OAI21X1_290/Y gnd vdd DFFPOSX1
XDFFPOSX1_2 OR2X2_1/B CLKBUF1_5/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XINVX1_372 AND2X2_3/Y gnd INVX1_372/Y vdd INVX1
XOAI21X1_551 BUFX2_10/Y INVX1_624/Y INVX1_623/Y gnd OAI21X1_551/Y vdd OAI21X1
XBUFX2_25 BUFX2_22/A gnd BUFX2_25/Y vdd BUFX2
XAOI22X1_99 AOI22X1_99/A AND2X2_77/Y AOI22X1_99/C AOI22X1_99/D gnd AOI22X1_99/Y vdd
+ AOI22X1
XDFFPOSX1_88 AND2X2_43/B CLKBUF1_24/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XOAI21X1_70 INVX1_67/Y AOI22X1_22/Y AOI22X1_23/Y gnd OAI21X1_70/Y vdd OAI21X1
XNAND2X1_85 AND2X2_1/B INVX1_64/A gnd NAND2X1_86/B vdd NAND2X1
XDFFPOSX1_154 AOI22X1_77/C CLKBUF1_37/Y OAI21X1_234/Y gnd vdd DFFPOSX1
XOAI21X1_515 INVX1_554/A INVX1_582/Y INVX1_581/Y gnd OAI21X1_516/C vdd OAI21X1
XAOI22X1_156 INVX1_532/A INVX1_531/Y INVX1_533/Y NAND2X1_458/Y gnd OAI21X1_478/B vdd
+ AOI22X1
XINVX1_336 INVX1_336/A gnd INVX1_336/Y vdd INVX1
XBUFX2_3 CLK gnd BUFX2_3/Y vdd BUFX2
XAOI22X1_63 AOI22X1_63/A AND2X2_56/Y AOI22X1_63/C NOR2X1_79/Y gnd AOI22X1_63/Y vdd
+ AOI22X1
XFILL_26_2_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XDFFPOSX1_118 AOI22X1_59/C CLKBUF1_16/Y OAI21X1_179/Y gnd vdd DFFPOSX1
XFILL_6_3_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XNAND2X1_49 OR2X2_4/B NOR2X1_21/Y gnd NAND2X1_49/Y vdd NAND2X1
XOAI21X1_34 INVX1_37/Y NOR2X1_21/Y NAND2X1_51/Y gnd OAI21X1_34/Y vdd OAI21X1
XDFFPOSX1_52 INVX1_72/A CLKBUF1_26/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XAOI22X1_120 INVX1_406/A INVX1_405/Y INVX1_407/Y NAND2X1_359/Y gnd OAI21X1_370/B vdd
+ AOI22X1
XOAI21X1_479 BUFX2_64/Y INVX1_540/Y INVX1_539/Y gnd OAI21X1_479/Y vdd OAI21X1
XINVX1_300 BUFX2_52/Y gnd INVX1_300/Y vdd INVX1
XNAND2X1_13 INVX1_476/A INVX1_296/A gnd NOR2X1_7/A vdd NAND2X1
XAOI22X1_27 AOI22X1_27/A AND2X2_35/Y AOI22X1_27/C NOR2X1_40/Y gnd AOI22X1_27/Y vdd
+ AOI22X1
XDFFPOSX1_16 INVX1_12/A CLKBUF1_5/Y NAND2X1_42/Y gnd vdd DFFPOSX1
XINVX1_264 BUFX2_32/Y gnd INVX1_264/Y vdd INVX1
XOAI21X1_443 BUFX2_130/Y INVX1_498/Y INVX1_497/Y gnd OAI21X1_444/C vdd OAI21X1
XNAND3X1_90 INVX1_575/A INVX1_288/Y INVX1_289/Y gnd NAND3X1_90/Y vdd NAND3X1
XINVX1_228 OR2X2_4/B gnd INVX1_228/Y vdd INVX1
XOAI21X1_407 BUFX2_114/Y INVX1_456/Y INVX1_455/Y gnd OAI21X1_407/Y vdd OAI21X1
XNAND3X1_54 INVX1_160/A INVX1_162/Y INVX1_163/Y gnd NAND3X1_54/Y vdd NAND3X1
XNAND2X1_521 INVX1_611/A NAND2X1_520/Y gnd NAND2X1_521/Y vdd NAND2X1
XNAND2X1_2 INVX1_588/A NAND2X1_2/B gnd NOR2X1_1/B vdd NAND2X1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_192 INVX1_375/A gnd INVX1_192/Y vdd INVX1
XOAI21X1_371 BUFX2_40/Y INVX1_414/Y INVX1_413/Y gnd OAI21X1_371/Y vdd OAI21X1
XAND2X2_123 INVX1_564/A INVX1_557/A gnd NOR2X1_210/B vdd AND2X2
XNAND3X1_18 INVX1_38/Y NAND2X1_61/Y OR2X2_4/Y gnd AND2X2_26/A vdd NAND3X1
XNAND2X1_485 AND2X2_42/A INVX1_566/Y gnd OAI21X1_507/B vdd NAND2X1
XAND2X2_96 AND2X2_96/A INVX1_431/A gnd AND2X2_96/Y vdd AND2X2
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XOAI21X1_335 INVX1_370/A INVX1_372/Y INVX1_371/Y gnd OAI21X1_336/C vdd OAI21X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XNAND2X1_449 INVX1_518/A BUFX2_65/Y gnd NAND2X1_450/B vdd NAND2X1
XAND2X2_60 BUFX2_16/Y AND2X2_60/B gnd AND2X2_60/Y vdd AND2X2
XINVX1_120 BUFX2_105/Y gnd NOR2X1_53/B vdd INVX1
XOAI21X1_299 INVX1_624/A INVX1_330/Y INVX1_329/Y gnd OAI21X1_300/C vdd OAI21X1
XNAND2X1_413 INVX1_475/A INVX1_478/A gnd NAND2X1_413/Y vdd NAND2X1
XAND2X2_24 OR2X2_2/A AND2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XNOR2X1_99 NOR2X1_99/A NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XOAI21X1_263 BUFX2_57/Y INVX1_286/Y OAI21X1_263/C gnd NAND3X1_91/C vdd OAI21X1
XNAND2X1_377 BUFX2_87/Y INVX1_429/Y gnd NAND2X1_377/Y vdd NAND2X1
XINVX1_625 AND2X2_21/A gnd INVX1_625/Y vdd INVX1
XNOR2X1_63 gnd INVX1_152/Y gnd NOR2X1_63/Y vdd NOR2X1
XOAI21X1_227 INVX1_244/Y INVX1_247/Y AOI22X1_75/C gnd OAI21X1_228/C vdd OAI21X1
XNAND2X1_341 INVX1_380/A NAND2X1_340/Y gnd NAND2X1_341/Y vdd NAND2X1
XCLKBUF1_51 BUFX2_4/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XINVX1_589 BUFX2_12/Y gnd INVX1_589/Y vdd INVX1
XNAND3X1_173 NOR2X1_223/Y NAND3X1_172/Y NAND3X1_173/C gnd NAND3X1_173/Y vdd NAND3X1
XFILL_22_1 gnd vdd FILL
XNOR2X1_27 NOR2X1_26/Y NOR2X1_27/B gnd NOR2X1_27/Y vdd NOR2X1
XOAI21X1_191 INVX1_206/Y OAI21X1_191/B OAI21X1_191/C gnd OAI21X1_191/Y vdd OAI21X1
XFILL_14_0_1 gnd vdd FILL
XNOR2X1_224 INVX1_574/A INVX1_575/Y gnd NOR2X1_224/Y vdd NOR2X1
XFILL_12_2_2 gnd vdd FILL
XNAND2X1_305 BUFX2_117/Y INVX1_335/Y gnd NAND2X1_305/Y vdd NAND2X1
XCLKBUF1_15 BUFX2_1/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XNAND3X1_137 NOR2X1_169/Y NAND3X1_136/Y NAND3X1_137/C gnd NAND3X1_137/Y vdd NAND3X1
XINVX1_553 INVX1_553/A gnd INVX1_553/Y vdd INVX1
XBUFX2_138 BUFX2_138/A gnd response_get[1] vdd BUFX2
XOAI21X1_155 INVX1_161/Y OAI21X1_155/B NOR2X1_65/Y gnd AOI21X1_24/C vdd OAI21X1
XNOR2X1_188 INVX1_490/A INVX1_491/Y gnd NOR2X1_188/Y vdd NOR2X1
XNAND2X1_269 INVX1_293/A INVX1_296/A gnd OAI21X1_271/B vdd NAND2X1
XDFFPOSX1_335 INVX1_122/A CLKBUF1_36/Y OAI21X1_508/Y gnd vdd DFFPOSX1
XBUFX2_102 BUFX2_98/A gnd INVX1_601/A vdd BUFX2
XINVX1_517 BUFX2_93/Y gnd INVX1_517/Y vdd INVX1
XNAND3X1_101 NOR2X1_115/Y NAND3X1_100/Y OAI21X1_294/Y gnd NAND3X1_101/Y vdd NAND3X1
XXNOR2X1_62 INVX1_463/A BUFX2_83/Y gnd XNOR2X1_62/Y vdd XNOR2X1
XOAI21X1_119 INVX1_123/Y AOI22X1_38/Y AOI22X1_39/Y gnd DFFPOSX1_79/D vdd OAI21X1
XNOR2X1_152 INVX1_406/A INVX1_407/Y gnd NOR2X1_152/Y vdd NOR2X1
XNAND2X1_233 INVX1_282/A INVX1_275/A gnd NOR2X1_93/A vdd NAND2X1
XINVX1_481 BUFX2_34/Y gnd INVX1_481/Y vdd INVX1
XFILL_13_3_0 gnd vdd FILL
XDFFPOSX1_299 INVX1_508/A CLKBUF1_12/Y OAI21X1_454/Y gnd vdd DFFPOSX1
XXNOR2X1_26 BUFX2_92/Y INVX1_209/A gnd XNOR2X1_26/Y vdd XNOR2X1
XNOR2X1_116 AND2X2_18/B INVX1_323/Y gnd AOI22X1_97/D vdd NOR2X1
XNAND2X1_197 AND2X2_10/B INVX1_204/A gnd NAND2X1_198/B vdd NAND2X1
XINVX1_445 INVX1_157/A gnd INVX1_445/Y vdd INVX1
XDFFPOSX1_263 INVX1_157/A CLKBUF1_15/Y OAI21X1_400/Y gnd vdd DFFPOSX1
XFILL_21_0_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XBUFX2_98 BUFX2_98/A gnd BUFX2_98/Y vdd BUFX2
XFILL_19_2_2 gnd vdd FILL
XNAND2X1_161 BUFX2_48/Y INVX1_160/Y gnd OAI21X1_155/B vdd NAND2X1
XAOI21X1_59 INVX1_408/Y AOI21X1_59/B AOI21X1_59/C gnd AOI21X1_59/Y vdd AOI21X1
XDFFPOSX1_227 AND2X2_88/B CLKBUF1_1/Y OAI21X1_346/Y gnd vdd DFFPOSX1
XINVX1_409 INVX1_409/A gnd INVX1_409/Y vdd INVX1
XBUFX2_62 BUFX2_65/A gnd BUFX2_62/Y vdd BUFX2
XNAND2X1_125 INVX1_114/A NAND2X1_124/Y gnd AOI22X1_37/A vdd NAND2X1
XINVX1_373 AND2X2_3/A gnd INVX1_373/Y vdd INVX1
XAOI21X1_23 INVX1_156/Y AOI21X1_23/B AOI21X1_23/C gnd AOI21X1_23/Y vdd AOI21X1
XDFFPOSX1_3 INVX1_16/A CLKBUF1_5/Y NAND3X1_13/Y gnd vdd DFFPOSX1
XOAI21X1_552 INVX1_624/A INVX1_622/Y OAI21X1_551/Y gnd OAI21X1_552/Y vdd OAI21X1
XDFFPOSX1_191 INVX1_319/A CLKBUF1_48/Y OAI21X1_292/Y gnd vdd DFFPOSX1
XBUFX2_26 BUFX2_22/A gnd BUFX2_26/Y vdd BUFX2
XFILL_20_3_0 gnd vdd FILL
XDFFPOSX1_155 INVX1_437/A CLKBUF1_29/Y OAI21X1_236/Y gnd vdd DFFPOSX1
XOAI21X1_71 INVX1_69/A INVX1_71/Y INVX1_70/Y gnd OAI21X1_72/C vdd OAI21X1
XDFFPOSX1_89 INVX1_133/A CLKBUF1_2/Y NAND3X1_47/Y gnd vdd DFFPOSX1
XNAND2X1_86 INVX1_65/A NAND2X1_86/B gnd AOI22X1_23/A vdd NAND2X1
XOAI21X1_516 INVX1_582/A INVX1_580/Y OAI21X1_516/C gnd NAND3X1_175/C vdd OAI21X1
XAOI22X1_157 NAND2X1_460/Y AND2X2_121/Y OAI21X1_475/C NOR2X1_206/Y gnd OAI21X1_478/C
+ vdd AOI22X1
XINVX1_337 BUFX2_117/Y gnd INVX1_337/Y vdd INVX1
XBUFX2_4 CLK gnd BUFX2_4/Y vdd BUFX2
XNAND2X1_50 INVX1_39/A NOR2X1_21/Y gnd OAI21X1_33/C vdd NAND2X1
XFILL_26_2_2 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XAOI22X1_64 INVX1_210/A INVX1_209/Y INVX1_211/Y AOI22X1_64/D gnd AOI22X1_64/Y vdd
+ AOI22X1
XDFFPOSX1_119 INVX1_193/A CLKBUF1_49/Y OAI21X1_181/Y gnd vdd DFFPOSX1
XAOI22X1_121 NAND2X1_361/Y AND2X2_94/Y AOI22X1_121/C NOR2X1_152/Y gnd AOI22X1_121/Y
+ vdd AOI22X1
XFILL_6_3_2 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XOAI21X1_35 INVX1_28/Y AND2X2_24/B NOR2X1_20/Y gnd AOI21X1_3/C vdd OAI21X1
XDFFPOSX1_53 INVX1_70/A CLKBUF1_26/Y NAND3X1_29/Y gnd vdd DFFPOSX1
XOAI21X1_480 INVX1_279/A INVX1_538/Y OAI21X1_479/Y gnd NAND3X1_163/C vdd OAI21X1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XAOI22X1_28 INVX1_84/A INVX1_83/Y INVX1_85/Y AOI22X1_28/D gnd OAI21X1_88/B vdd AOI22X1
XNAND2X1_14 INVX1_602/A INVX1_560/A gnd NOR2X1_7/B vdd NAND2X1
XDFFPOSX1_17 INVX1_13/A CLKBUF1_18/Y NAND2X1_43/Y gnd vdd DFFPOSX1
XOAI21X1_444 INVX1_498/A INVX1_496/Y OAI21X1_444/C gnd NAND3X1_151/C vdd OAI21X1
XINVX1_265 BUFX2_59/Y gnd INVX1_265/Y vdd INVX1
XNAND3X1_91 NOR2X1_104/Y NAND3X1_90/Y NAND3X1_91/C gnd NAND3X1_91/Y vdd NAND3X1
XFILL_27_3_0 gnd vdd FILL
XINVX1_229 BUFX2_34/Y gnd NOR2X1_87/B vdd INVX1
XOAI21X1_408 AND2X2_9/Y INVX1_454/Y OAI21X1_407/Y gnd OAI21X1_408/Y vdd OAI21X1
XNAND3X1_55 NOR2X1_65/Y NAND3X1_54/Y NAND3X1_55/C gnd NAND3X1_55/Y vdd NAND3X1
XNAND2X1_522 BUFX2_8/Y AND2X2_20/A gnd NAND2X1_522/Y vdd NAND2X1
XNAND2X1_3 INVX1_343/A INVX1_86/A gnd NOR2X1_2/A vdd NAND2X1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XINVX1_75 BUFX2_32/Y gnd INVX1_75/Y vdd INVX1
XOAI21X1_372 AND2X2_6/Y INVX1_412/Y OAI21X1_371/Y gnd OAI21X1_372/Y vdd OAI21X1
XNAND2X1_486 INVX1_566/A INVX1_569/Y gnd NAND2X1_486/Y vdd NAND2X1
XAND2X2_124 INVX1_564/A INVX1_550/A gnd AND2X2_124/Y vdd AND2X2
XNAND3X1_19 INVX1_39/A NAND3X1_19/B OR2X2_5/Y gnd NAND3X1_19/Y vdd NAND3X1
XAND2X2_97 AND2X2_96/A AND2X2_98/B gnd AND2X2_97/Y vdd AND2X2
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XOAI21X1_336 AND2X2_3/Y INVX1_370/Y OAI21X1_336/C gnd NAND3X1_115/C vdd OAI21X1
XNAND2X1_450 INVX1_520/A NAND2X1_450/B gnd NAND2X1_450/Y vdd NAND2X1
XAND2X2_61 AND2X2_6/Y INVX1_417/A gnd AND2X2_61/Y vdd AND2X2
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XOAI21X1_300 BUFX2_20/Y INVX1_328/Y OAI21X1_300/C gnd NAND3X1_103/C vdd OAI21X1
XNAND2X1_414 BUFX2_133/Y INVX1_475/Y gnd NAND2X1_414/Y vdd NAND2X1
XAND2X2_25 OR2X2_4/A OR2X2_4/B gnd AND2X2_25/Y vdd AND2X2
XOAI21X1_264 INVX1_286/Y INVX1_289/Y AOI22X1_87/C gnd OAI21X1_265/C vdd OAI21X1
XNAND2X1_378 INVX1_427/A BUFX2_116/Y gnd NAND2X1_379/B vdd NAND2X1
XNOR2X1_64 AND2X2_7/B INVX1_155/Y gnd NOR2X1_64/Y vdd NOR2X1
XINVX1_626 INVX1_626/A gnd INVX1_626/Y vdd INVX1
XOAI21X1_228 INVX1_248/Y NAND2X1_228/Y OAI21X1_228/C gnd OAI21X1_228/Y vdd OAI21X1
XNAND2X1_342 BUFX2_79/Y INVX1_387/A gnd OAI21X1_350/B vdd NAND2X1
XNAND3X1_174 INVX1_580/A INVX1_582/Y INVX1_583/Y gnd NAND3X1_175/B vdd NAND3X1
XINVX1_590 INVX1_590/A gnd INVX1_590/Y vdd INVX1
XNOR2X1_28 NOR2X1_28/A NOR2X1_28/B gnd BUFX2_44/A vdd NOR2X1
XFILL_22_2 gnd vdd FILL
XOAI21X1_192 INVX1_203/Y NAND2X1_195/Y NOR2X1_78/Y gnd AOI21X1_30/C vdd OAI21X1
XFILL_14_0_2 gnd vdd FILL
XNOR2X1_225 gnd INVX1_579/Y gnd NOR2X1_225/Y vdd NOR2X1
XNAND2X1_306 BUFX2_22/Y INVX1_338/Y gnd NAND2X1_306/Y vdd NAND2X1
XCLKBUF1_16 BUFX2_5/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XBUFX2_139 BUFX2_139/A gnd response_get[2] vdd BUFX2
XNAND3X1_138 BUFX2_114/Y INVX1_456/Y INVX1_457/Y gnd NAND3X1_138/Y vdd NAND3X1
XINVX1_554 INVX1_554/A gnd INVX1_554/Y vdd INVX1
XOAI21X1_156 INVX1_165/Y AOI22X1_50/Y AOI22X1_51/Y gnd OAI21X1_156/Y vdd OAI21X1
XNOR2X1_189 gnd INVX1_495/Y gnd NOR2X1_189/Y vdd NOR2X1
XNAND2X1_270 BUFX2_100/Y INVX1_293/Y gnd OAI21X1_272/B vdd NAND2X1
XDFFPOSX1_336 AND2X2_16/A CLKBUF1_23/Y AOI21X1_82/Y gnd vdd DFFPOSX1
XBUFX2_103 BUFX2_103/A gnd INVX1_106/A vdd BUFX2
XNAND3X1_102 INVX1_624/A INVX1_330/Y INVX1_331/Y gnd NAND3X1_102/Y vdd NAND3X1
XINVX1_518 INVX1_518/A gnd INVX1_518/Y vdd INVX1
XNOR2X1_153 gnd INVX1_411/Y gnd NOR2X1_153/Y vdd NOR2X1
XXNOR2X1_63 BUFX2_132/Y BUFX2_91/Y gnd XNOR2X1_63/Y vdd XNOR2X1
XOAI21X1_120 INVX1_125/A NOR2X1_56/B INVX1_126/Y gnd OAI21X1_121/C vdd OAI21X1
XFILL_15_1_0 gnd vdd FILL
XNAND2X1_234 NOR2X1_99/A INVX1_289/A gnd NOR2X1_93/B vdd NAND2X1
XINVX1_482 BUFX2_134/Y gnd INVX1_482/Y vdd INVX1
XFILL_13_3_1 gnd vdd FILL
XDFFPOSX1_300 INVX1_506/A CLKBUF1_3/Y AOI21X1_73/Y gnd vdd DFFPOSX1
XXNOR2X1_27 INVX1_209/A BUFX2_55/Y gnd AOI21X1_32/B vdd XNOR2X1
XNAND2X1_198 INVX1_205/A NAND2X1_198/B gnd AOI22X1_63/A vdd NAND2X1
XNOR2X1_117 gnd INVX1_327/Y gnd NOR2X1_117/Y vdd NOR2X1
XDFFPOSX1_264 AND2X2_7/A CLKBUF1_10/Y AOI21X1_64/Y gnd vdd DFFPOSX1
XINVX1_446 BUFX2_31/Y gnd INVX1_446/Y vdd INVX1
XFILL_21_0_2 gnd vdd FILL
XFILL_1_1_2 gnd vdd FILL
XBUFX2_99 BUFX2_98/A gnd BUFX2_99/Y vdd BUFX2
XNAND2X1_162 INVX1_160/A INVX1_163/Y gnd AOI22X1_50/D vdd NAND2X1
XXOR2X1_1 OR2X2_5/A OR2X2_3/B gnd XOR2X1_1/Y vdd XOR2X1
XINVX1_410 AND2X2_47/B gnd INVX1_410/Y vdd INVX1
XAOI21X1_60 INVX1_415/Y AOI21X1_60/B AOI21X1_60/C gnd AOI21X1_60/Y vdd AOI21X1
XDFFPOSX1_228 INVX1_380/A CLKBUF1_19/Y AOI21X1_55/Y gnd vdd DFFPOSX1
XBUFX2_63 BUFX2_65/A gnd BUFX2_63/Y vdd BUFX2
XNAND2X1_126 AND2X2_42/A INVX1_121/A gnd OAI21X1_117/B vdd NAND2X1
XINVX1_374 AND2X2_86/B gnd INVX1_374/Y vdd INVX1
XAOI21X1_24 INVX1_163/Y XNOR2X1_19/Y AOI21X1_24/C gnd AOI21X1_24/Y vdd AOI21X1
XDFFPOSX1_4 INVX1_18/A CLKBUF1_18/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XOAI21X1_553 INVX1_622/Y INVX1_625/Y AOI22X1_183/C gnd OAI21X1_553/Y vdd OAI21X1
XDFFPOSX1_192 INVX1_317/A CLKBUF1_44/Y AOI21X1_46/Y gnd vdd DFFPOSX1
XBUFX2_27 RST_N gnd INVX1_96/A vdd BUFX2
XFILL_22_1_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XNAND2X1_87 INVX1_69/A INVX1_72/A gnd NAND2X1_87/Y vdd NAND2X1
XFILL_20_3_1 gnd vdd FILL
XDFFPOSX1_90 AOI22X1_45/C CLKBUF1_8/Y OAI21X1_135/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 INVX1_254/A CLKBUF1_37/Y AOI21X1_37/Y gnd vdd DFFPOSX1
XOAI21X1_72 BUFX2_43/Y INVX1_69/Y OAI21X1_72/C gnd OAI21X1_72/Y vdd OAI21X1
XBUFX2_5 CLK gnd BUFX2_5/Y vdd BUFX2
XAOI22X1_158 INVX1_539/A INVX1_538/Y INVX1_540/Y NAND2X1_463/Y gnd OAI21X1_484/B vdd
+ AOI22X1
XINVX1_338 INVX1_338/A gnd INVX1_338/Y vdd INVX1
XOAI21X1_517 INVX1_580/Y INVX1_583/Y OAI21X1_517/C gnd OAI21X1_518/C vdd OAI21X1
XFILL_28_0_2 gnd vdd FILL
XFILL_8_1_2 gnd vdd FILL
XNAND2X1_51 INVX1_38/A NOR2X1_21/Y gnd NAND2X1_51/Y vdd NAND2X1
XOAI21X1_36 NOR2X1_22/Y AOI21X1_4/Y BUFX2_137/A gnd NAND2X1_53/A vdd OAI21X1
XAOI22X1_65 AOI22X1_65/A AND2X2_58/Y AOI22X1_65/C NOR2X1_82/Y gnd AOI22X1_65/Y vdd
+ AOI22X1
XDFFPOSX1_120 INVX1_191/A CLKBUF1_49/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XAOI22X1_122 INVX1_413/A INVX1_412/Y INVX1_414/Y NAND2X1_364/Y gnd OAI21X1_376/B vdd
+ AOI22X1
XOAI21X1_481 INVX1_538/Y INVX1_541/Y AOI22X1_159/C gnd OAI21X1_482/C vdd OAI21X1
XDFFPOSX1_54 AOI22X1_27/C CLKBUF1_51/Y OAI21X1_80/Y gnd vdd DFFPOSX1
XINVX1_302 INVX1_293/A gnd INVX1_302/Y vdd INVX1
XAOI22X1_29 AOI22X1_29/A AND2X2_37/Y OAI21X1_85/C NOR2X1_43/Y gnd OAI21X1_88/C vdd
+ AOI22X1
XDFFPOSX1_18 OR2X2_2/B CLKBUF1_28/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XNAND2X1_15 INVX1_133/A INVX1_91/A gnd NOR2X1_8/A vdd NAND2X1
XOAI21X1_445 INVX1_496/Y INVX1_499/Y OAI21X1_445/C gnd OAI21X1_445/Y vdd OAI21X1
XINVX1_266 NOR2X1_99/A gnd INVX1_266/Y vdd INVX1
XFILL_13_1 gnd vdd FILL
XNAND3X1_92 INVX1_293/A INVX1_295/Y INVX1_296/Y gnd NAND3X1_92/Y vdd NAND3X1
XFILL_27_3_1 gnd vdd FILL
XNAND3X1_56 INVX1_167/A INVX1_169/Y INVX1_170/Y gnd NAND3X1_56/Y vdd NAND3X1
XINVX1_230 AND2X2_6/Y gnd INVX1_230/Y vdd INVX1
XOAI21X1_409 INVX1_454/Y INVX1_457/Y OAI21X1_409/C gnd OAI21X1_410/C vdd OAI21X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_523 INVX1_160/A INVX1_615/Y gnd OAI21X1_549/B vdd NAND2X1
XNAND2X1_4 NAND2X1_4/A INVX1_378/A gnd NOR2X1_2/B vdd NAND2X1
XINVX1_194 BUFX2_31/Y gnd INVX1_194/Y vdd INVX1
XOAI21X1_373 INVX1_412/Y INVX1_415/Y OAI21X1_373/C gnd OAI21X1_374/C vdd OAI21X1
XAND2X2_125 INVX1_557/A INVX1_550/A gnd AND2X2_125/Y vdd AND2X2
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XNAND2X1_487 INVX1_567/A AND2X2_42/A gnd NAND2X1_488/B vdd NAND2X1
XNAND3X1_20 INVX1_41/A INVX1_43/Y INVX1_44/Y gnd NAND3X1_21/B vdd NAND3X1
XAND2X2_98 INVX1_431/A AND2X2_98/B gnd AND2X2_98/Y vdd AND2X2
XINVX1_40 INVX1_89/A gnd INVX1_40/Y vdd INVX1
XOAI21X1_337 INVX1_370/Y INVX1_373/Y OAI21X1_337/C gnd OAI21X1_338/C vdd OAI21X1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XNAND2X1_451 BUFX2_63/Y AND2X2_13/A gnd NAND2X1_451/Y vdd NAND2X1
XAND2X2_62 INVX1_237/A INVX1_241/A gnd AND2X2_62/Y vdd AND2X2
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XNAND2X1_415 INVX1_475/A INVX1_478/Y gnd AOI22X1_140/D vdd NAND2X1
XOAI21X1_301 INVX1_328/Y INVX1_331/Y AOI22X1_99/C gnd OAI21X1_302/C vdd OAI21X1
XAND2X2_26 AND2X2_26/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XOAI21X1_265 INVX1_290/Y OAI21X1_265/B OAI21X1_265/C gnd OAI21X1_265/Y vdd OAI21X1
XNAND2X1_379 INVX1_429/A NAND2X1_379/B gnd NAND2X1_379/Y vdd NAND2X1
XNOR2X1_65 gnd NOR2X1_65/B gnd NOR2X1_65/Y vdd NOR2X1
XINVX1_627 INVX1_627/A gnd INVX1_627/Y vdd INVX1
XOAI21X1_229 INVX1_245/Y OAI21X1_229/B NOR2X1_91/Y gnd AOI21X1_36/C vdd OAI21X1
XNAND2X1_343 BUFX2_37/Y INVX1_384/Y gnd OAI21X1_351/B vdd NAND2X1
XNAND3X1_175 NOR2X1_225/Y NAND3X1_175/B NAND3X1_175/C gnd NAND3X1_175/Y vdd NAND3X1
XINVX1_591 INVX1_46/A gnd INVX1_591/Y vdd INVX1
XOAI21X1_193 INVX1_207/Y AOI22X1_62/Y AOI22X1_63/Y gnd OAI21X1_193/Y vdd OAI21X1
XNOR2X1_29 gnd INVX1_40/Y gnd NOR2X1_29/Y vdd NOR2X1
XNAND2X1_307 INVX1_336/A BUFX2_117/Y gnd NAND2X1_307/Y vdd NAND2X1
XNOR2X1_226 INVX1_581/A INVX1_582/Y gnd NOR2X1_226/Y vdd NOR2X1
XNAND3X1_139 NOR2X1_171/Y NAND3X1_138/Y OAI21X1_408/Y gnd NAND3X1_139/Y vdd NAND3X1
XCLKBUF1_17 BUFX2_2/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XINVX1_555 INVX1_555/A gnd INVX1_555/Y vdd INVX1
XBUFX2_140 BUFX2_140/A gnd response_get[3] vdd BUFX2
XOAI21X1_157 INVX1_167/A INVX1_169/Y INVX1_168/Y gnd OAI21X1_157/Y vdd OAI21X1
XNOR2X1_190 INVX1_497/A INVX1_498/Y gnd NOR2X1_190/Y vdd NOR2X1
XNAND2X1_271 INVX1_293/A INVX1_296/Y gnd AOI22X1_88/D vdd NAND2X1
XDFFPOSX1_337 INVX1_567/A CLKBUF1_36/Y NAND3X1_171/Y gnd vdd DFFPOSX1
XNAND3X1_103 NOR2X1_117/Y NAND3X1_102/Y NAND3X1_103/C gnd NAND3X1_103/Y vdd NAND3X1
XINVX1_519 BUFX2_65/Y gnd INVX1_519/Y vdd INVX1
XBUFX2_104 BUFX2_103/A gnd INVX1_97/A vdd BUFX2
XNOR2X1_154 INVX1_413/A INVX1_414/Y gnd NOR2X1_154/Y vdd NOR2X1
XXNOR2X1_64 BUFX2_133/Y BUFX2_98/Y gnd XNOR2X1_64/Y vdd XNOR2X1
XOAI21X1_121 BUFX2_82/Y INVX1_125/Y OAI21X1_121/C gnd NAND3X1_45/C vdd OAI21X1
XNAND2X1_235 INVX1_251/A INVX1_254/A gnd NAND2X1_235/Y vdd NAND2X1
XFILL_15_1_1 gnd vdd FILL
XINVX1_483 INVX1_483/A gnd INVX1_483/Y vdd INVX1
XFILL_13_3_2 gnd vdd FILL
XDFFPOSX1_301 NAND2X1_2/B CLKBUF1_12/Y NAND3X1_153/Y gnd vdd DFFPOSX1
XXNOR2X1_28 BUFX2_67/Y BUFX2_16/Y gnd XNOR2X1_28/Y vdd XNOR2X1
XNAND2X1_199 INVX1_240/A INVX1_233/A gnd NOR2X1_80/A vdd NAND2X1
XNOR2X1_118 AND2X2_21/B INVX1_330/Y gnd AOI22X1_99/D vdd NOR2X1
XDFFPOSX1_265 INVX1_441/A CLKBUF1_10/Y NAND3X1_135/Y gnd vdd DFFPOSX1
XINVX1_447 BUFX2_113/Y gnd INVX1_447/Y vdd INVX1
XNAND2X1_163 INVX1_161/A BUFX2_48/Y gnd NAND2X1_163/Y vdd NAND2X1
XINVX1_411 BUFX2_28/Y gnd INVX1_411/Y vdd INVX1
XAOI21X1_61 INVX1_422/Y XNOR2X1_56/Y AOI21X1_61/C gnd AOI21X1_61/Y vdd AOI21X1
XDFFPOSX1_229 INVX1_378/A CLKBUF1_1/Y NAND3X1_117/Y gnd vdd DFFPOSX1
XBUFX2_64 BUFX2_65/A gnd BUFX2_64/Y vdd BUFX2
XNAND2X1_127 BUFX2_105/Y INVX1_118/Y gnd OAI21X1_118/B vdd NAND2X1
XDFFPOSX1_5 INVX1_20/A CLKBUF1_12/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XDFFPOSX1_193 AND2X2_12/B CLKBUF1_40/Y NAND3X1_99/Y gnd vdd DFFPOSX1
XAOI21X1_25 INVX1_170/Y AOI21X1_25/B AOI21X1_25/C gnd AOI21X1_25/Y vdd AOI21X1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XOAI21X1_554 INVX1_626/Y NAND2X1_527/Y OAI21X1_553/Y gnd OAI21X1_554/Y vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XBUFX2_28 RST_N gnd BUFX2_28/Y vdd BUFX2
XFILL_22_1_1 gnd vdd FILL
XFILL_20_3_2 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XNAND2X1_88 BUFX2_43/Y INVX1_69/Y gnd OAI21X1_75/B vdd NAND2X1
XDFFPOSX1_91 OR2X2_3/B CLKBUF1_8/Y OAI21X1_137/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 NOR2X1_95/A CLKBUF1_13/Y NAND3X1_81/Y gnd vdd DFFPOSX1
XAOI22X1_159 NAND2X1_465/Y AND2X2_122/Y AOI22X1_159/C NOR2X1_208/Y gnd OAI21X1_484/C
+ vdd AOI22X1
XOAI21X1_73 INVX1_69/Y INVX1_72/Y AOI22X1_25/C gnd OAI21X1_73/Y vdd OAI21X1
XBUFX2_6 CLK gnd BUFX2_6/Y vdd BUFX2
XINVX1_339 INVX1_46/A gnd INVX1_339/Y vdd INVX1
XOAI21X1_518 INVX1_584/Y OAI21X1_518/B OAI21X1_518/C gnd OAI21X1_518/Y vdd OAI21X1
XAOI22X1_66 INVX1_217/A INVX1_216/Y INVX1_218/Y AOI22X1_66/D gnd AOI22X1_66/Y vdd
+ AOI22X1
XOAI21X1_37 INVX1_27/Y OR2X2_2/B OAI21X1_37/C gnd AOI22X1_9/D vdd OAI21X1
XNAND2X1_52 EN_response_get INVX1_27/Y gnd AND2X2_24/B vdd NAND2X1
XDFFPOSX1_55 INVX1_81/A CLKBUF1_26/Y OAI21X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 AND2X2_3/B CLKBUF1_16/Y NAND3X1_63/Y gnd vdd DFFPOSX1
XAOI22X1_123 AOI22X1_123/A AND2X2_95/Y OAI21X1_373/C NOR2X1_154/Y gnd OAI21X1_376/C
+ vdd AOI22X1
XINVX1_303 AND2X2_71/B gnd INVX1_303/Y vdd INVX1
XOAI21X1_482 INVX1_542/Y OAI21X1_482/B OAI21X1_482/C gnd OAI21X1_482/Y vdd OAI21X1
XAOI22X1_30 INVX1_91/A INVX1_90/Y INVX1_92/Y AOI22X1_30/D gnd OAI21X1_94/B vdd AOI22X1
XDFFPOSX1_19 INVX1_28/A CLKBUF1_28/Y NAND3X1_15/Y gnd vdd DFFPOSX1
XNAND2X1_16 INVX1_217/A NOR2X1_71/A gnd NOR2X1_8/B vdd NAND2X1
XOAI21X1_446 INVX1_500/Y OAI21X1_446/B OAI21X1_445/Y gnd OAI21X1_446/Y vdd OAI21X1
XINVX1_267 BUFX2_68/Y gnd NOR2X1_99/B vdd INVX1
XFILL_13_2 gnd vdd FILL
XNAND3X1_93 NAND3X1_93/A NAND3X1_92/Y NAND3X1_93/C gnd NAND3X1_93/Y vdd NAND3X1
XINVX1_231 AND2X2_6/B gnd INVX1_231/Y vdd INVX1
XFILL_9_2_1 gnd vdd FILL
XFILL_27_3_2 gnd vdd FILL
XNAND3X1_57 NOR2X1_68/Y NAND3X1_56/Y NAND3X1_57/C gnd NAND3X1_57/Y vdd NAND3X1
XOAI21X1_410 INVX1_458/Y OAI21X1_410/B OAI21X1_410/C gnd OAI21X1_410/Y vdd OAI21X1
XNAND2X1_524 BUFX2_8/Y INVX1_618/Y gnd AOI22X1_180/D vdd NAND2X1
XNAND2X1_5 INVX1_385/A NAND2X1_5/B gnd NOR2X1_3/A vdd NAND2X1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_195 AND2X2_8/Y gnd INVX1_195/Y vdd INVX1
XOAI21X1_374 INVX1_416/Y OAI21X1_374/B OAI21X1_374/C gnd OAI21X1_374/Y vdd OAI21X1
XAND2X2_126 BUFX2_75/Y INVX1_88/A gnd AND2X2_126/Y vdd AND2X2
XNAND2X1_488 AND2X2_16/A NAND2X1_488/B gnd AOI22X1_167/A vdd NAND2X1
XNAND3X1_21 NOR2X1_29/Y NAND3X1_21/B OAI21X1_47/Y gnd NAND3X1_21/Y vdd NAND3X1
XAND2X2_99 BUFX2_79/Y AND2X2_99/B gnd AND2X2_99/Y vdd AND2X2
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XOAI21X1_338 INVX1_374/Y NAND2X1_329/Y OAI21X1_338/C gnd OAI21X1_338/Y vdd OAI21X1
XINVX1_159 BUFX2_35/Y gnd NOR2X1_65/B vdd INVX1
XNAND2X1_452 INVX1_69/A INVX1_524/Y gnd OAI21X1_471/B vdd NAND2X1
XAND2X2_63 INVX1_244/A AND2X2_63/B gnd AND2X2_63/Y vdd AND2X2
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XOAI21X1_302 INVX1_332/Y NAND2X1_296/Y OAI21X1_302/C gnd OAI21X1_302/Y vdd OAI21X1
XNAND2X1_416 INVX1_476/A BUFX2_133/Y gnd NAND2X1_417/B vdd NAND2X1
XAND2X2_27 OR2X2_5/A OR2X2_4/B gnd AND2X2_27/Y vdd AND2X2
XOAI21X1_266 INVX1_287/Y NAND2X1_263/Y NOR2X1_104/Y gnd AOI21X1_42/C vdd OAI21X1
XNAND2X1_380 BUFX2_97/Y INVX1_436/A gnd NAND2X1_380/Y vdd NAND2X1
XNOR2X1_66 INVX1_161/A INVX1_162/Y gnd NOR2X1_66/Y vdd NOR2X1
XOAI21X1_230 INVX1_249/Y AOI22X1_74/Y AOI22X1_75/Y gnd OAI21X1_230/Y vdd OAI21X1
XNAND2X1_344 BUFX2_81/Y INVX1_387/Y gnd AOI22X1_114/D vdd NAND2X1
XNAND3X1_176 BUFX2_24/Y INVX1_589/Y INVX1_590/Y gnd NAND3X1_176/Y vdd NAND3X1
XINVX1_592 INVX1_592/A gnd INVX1_592/Y vdd INVX1
XNOR2X1_30 INVX1_42/A INVX1_43/Y gnd NOR2X1_30/Y vdd NOR2X1
XOAI21X1_194 INVX1_209/A INVX1_211/Y INVX1_210/Y gnd OAI21X1_195/C vdd OAI21X1
XNAND2X1_308 INVX1_338/A NAND2X1_307/Y gnd AOI22X1_101/A vdd NAND2X1
XNOR2X1_227 INVX1_606/A INVX1_599/A gnd NOR2X1_227/Y vdd NOR2X1
XNAND3X1_140 BUFX2_83/Y INVX1_463/Y INVX1_464/Y gnd NAND3X1_140/Y vdd NAND3X1
XBUFX2_141 BUFX2_141/A gnd response_get[4] vdd BUFX2
XINVX1_556 INVX1_437/A gnd INVX1_556/Y vdd INVX1
XCLKBUF1_18 BUFX2_4/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XOAI21X1_158 BUFX2_85/Y INVX1_167/Y OAI21X1_157/Y gnd NAND3X1_57/C vdd OAI21X1
XNOR2X1_191 INVX1_522/A INVX1_515/A gnd NOR2X1_191/Y vdd NOR2X1
XNAND2X1_272 INVX1_294/A BUFX2_100/Y gnd NAND2X1_273/B vdd NAND2X1
XBUFX2_105 BUFX2_103/A gnd BUFX2_105/Y vdd BUFX2
XINVX1_520 INVX1_520/A gnd INVX1_520/Y vdd INVX1
XNAND3X1_104 BUFX2_22/Y INVX1_337/Y INVX1_338/Y gnd NAND3X1_104/Y vdd NAND3X1
XDFFPOSX1_338 AOI22X1_169/C CLKBUF1_38/Y OAI21X1_512/Y gnd vdd DFFPOSX1
XXNOR2X1_65 INVX1_484/A BUFX2_134/Y gnd AOI21X1_70/B vdd XNOR2X1
XOAI21X1_122 INVX1_125/Y INVX1_128/Y AOI22X1_41/C gnd OAI21X1_123/C vdd OAI21X1
XNOR2X1_155 AND2X2_96/A INVX1_431/A gnd NOR2X1_156/A vdd NOR2X1
XNAND2X1_236 BUFX2_95/Y INVX1_251/Y gnd NAND2X1_236/Y vdd NAND2X1
XFILL_15_1_2 gnd vdd FILL
XDFFPOSX1_302 AOI22X1_151/C CLKBUF1_5/Y OAI21X1_458/Y gnd vdd DFFPOSX1
XINVX1_484 INVX1_484/A gnd INVX1_484/Y vdd INVX1
XXNOR2X1_29 BUFX2_14/Y AND2X2_6/Y gnd XNOR2X1_29/Y vdd XNOR2X1
XNAND2X1_200 INVX1_224/A INVX1_247/A gnd NOR2X1_80/B vdd NAND2X1
XNOR2X1_119 INVX1_354/A AND2X2_80/A gnd NOR2X1_119/Y vdd NOR2X1
XDFFPOSX1_266 AOI22X1_133/C CLKBUF1_45/Y OAI21X1_404/Y gnd vdd DFFPOSX1
XINVX1_448 INVX1_448/A gnd INVX1_448/Y vdd INVX1
XNAND2X1_164 INVX1_163/A NAND2X1_163/Y gnd AOI22X1_51/A vdd NAND2X1
XFILL_26_1 gnd vdd FILL
XAOI21X1_62 INVX1_429/Y AOI21X1_62/B AOI21X1_62/C gnd AOI21X1_62/Y vdd AOI21X1
XINVX1_412 BUFX2_40/Y gnd INVX1_412/Y vdd INVX1
XDFFPOSX1_230 OAI21X1_349/C CLKBUF1_41/Y OAI21X1_350/Y gnd vdd DFFPOSX1
XFILL_16_2_0 gnd vdd FILL
XBUFX2_65 BUFX2_65/A gnd BUFX2_65/Y vdd BUFX2
XNAND2X1_128 AND2X2_42/A INVX1_121/Y gnd AOI22X1_38/D vdd NAND2X1
XAOI21X1_26 INVX1_177/Y AOI21X1_26/B AOI21X1_26/C gnd AOI21X1_26/Y vdd AOI21X1
XDFFPOSX1_6 INVX1_21/A CLKBUF1_18/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_194 AOI22X1_97/C CLKBUF1_7/Y OAI21X1_296/Y gnd vdd DFFPOSX1
XINVX1_376 INVX1_96/A gnd INVX1_376/Y vdd INVX1
XOAI21X1_555 INVX1_623/Y NAND2X1_528/Y NOR2X1_243/Y gnd AOI21X1_90/C vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XBUFX2_29 RST_N gnd INVX1_89/A vdd BUFX2
XFILL_22_1_2 gnd vdd FILL
XFILL_2_2_2 gnd vdd FILL
XOAI21X1_74 INVX1_73/Y NAND2X1_87/Y OAI21X1_73/Y gnd OAI21X1_74/Y vdd OAI21X1
XNAND2X1_89 INVX1_69/A INVX1_72/Y gnd AOI22X1_24/D vdd NAND2X1
XDFFPOSX1_92 INVX1_142/A CLKBUF1_10/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XAOI22X1_160 NAND2X1_4/A INVX1_545/Y INVX1_547/Y AOI22X1_160/D gnd OAI21X1_490/B vdd
+ AOI22X1
XOAI21X1_519 INVX1_581/Y NAND2X1_495/Y NOR2X1_225/Y gnd AOI21X1_84/C vdd OAI21X1
XINVX1_340 AND2X2_79/B gnd INVX1_340/Y vdd INVX1
XDFFPOSX1_158 AOI22X1_79/C CLKBUF1_37/Y OAI21X1_240/Y gnd vdd DFFPOSX1
XBUFX2_7 CLK gnd BUFX2_7/Y vdd BUFX2
XAOI22X1_67 AOI22X1_67/A AND2X2_59/Y AOI22X1_67/C NOR2X1_84/Y gnd AOI22X1_67/Y vdd
+ AOI22X1
XDFFPOSX1_122 AOI22X1_61/C CLKBUF1_49/Y OAI21X1_185/Y gnd vdd DFFPOSX1
XOAI21X1_38 NOR2X1_22/Y AOI21X1_4/Y BUFX2_138/A gnd NAND2X1_54/A vdd OAI21X1
XNAND2X1_53 NAND2X1_53/A AOI22X1_8/Y gnd NAND2X1_53/Y vdd NAND2X1
XDFFPOSX1_56 INVX1_79/A CLKBUF1_51/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XAOI22X1_124 INVX1_420/A INVX1_419/Y INVX1_421/Y AOI22X1_124/D gnd OAI21X1_382/B vdd
+ AOI22X1
XOAI21X1_483 INVX1_539/Y NAND2X1_462/Y NOR2X1_207/Y gnd AOI21X1_78/C vdd OAI21X1
XINVX1_304 AND2X2_73/B gnd INVX1_304/Y vdd INVX1
XAOI22X1_31 AOI22X1_31/A AND2X2_38/Y AOI22X1_31/C NOR2X1_45/Y gnd OAI21X1_94/C vdd
+ AOI22X1
XFILL_23_2_0 gnd vdd FILL
XNAND2X1_17 INVX1_301/A NOR2X1_97/A gnd INVX1_1/A vdd NAND2X1
XFILL_3_3_0 gnd vdd FILL
XDFFPOSX1_20 INVX1_30/A CLKBUF1_20/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XOAI21X1_447 INVX1_497/Y NAND2X1_429/Y NOR2X1_189/Y gnd AOI21X1_72/C vdd OAI21X1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XNAND3X1_94 BUFX2_52/Y INVX1_302/Y INVX1_303/Y gnd NAND3X1_94/Y vdd NAND3X1
XFILL_13_3 gnd vdd FILL
XINVX1_232 BUFX2_14/Y gnd NOR2X1_88/B vdd INVX1
XFILL_9_2_2 gnd vdd FILL
XOAI21X1_411 INVX1_455/Y OAI21X1_411/B NOR2X1_171/Y gnd AOI21X1_66/C vdd OAI21X1
XNAND2X1_525 INVX1_616/A INVX1_160/A gnd NAND2X1_526/B vdd NAND2X1
XNAND3X1_58 BUFX2_54/Y NOR2X1_71/B INVX1_177/Y gnd NAND3X1_58/Y vdd NAND3X1
XNAND2X1_6 INVX1_420/A NAND2X1_6/B gnd NOR2X1_3/B vdd NAND2X1
XINVX1_78 BUFX2_42/Y gnd INVX1_78/Y vdd INVX1
XOAI21X1_375 INVX1_413/Y OAI21X1_375/B NOR2X1_153/Y gnd AOI21X1_60/C vdd OAI21X1
XINVX1_196 AND2X2_8/B gnd INVX1_196/Y vdd INVX1
XAND2X2_127 BUFX2_94/Y INVX1_437/A gnd AND2X2_127/Y vdd AND2X2
XNAND3X1_22 BUFX2_56/Y INVX1_50/Y INVX1_51/Y gnd NAND3X1_22/Y vdd NAND3X1
XNAND2X1_489 BUFX2_124/Y INVX1_576/A gnd OAI21X1_512/B vdd NAND2X1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XOAI21X1_339 INVX1_371/Y OAI21X1_339/B NOR2X1_135/Y gnd AOI21X1_54/C vdd OAI21X1
XNAND2X1_453 BUFX2_66/Y INVX1_527/Y gnd NAND2X1_453/Y vdd NAND2X1
XAND2X2_64 NOR2X1_95/A AND2X2_64/B gnd INVX1_251/A vdd AND2X2
XOAI21X1_303 INVX1_329/Y NAND2X1_297/Y NOR2X1_117/Y gnd AOI21X1_48/C vdd OAI21X1
XINVX1_124 INVX1_96/A gnd NOR2X1_55/B vdd INVX1
XNAND2X1_417 INVX1_478/A NAND2X1_417/B gnd NAND2X1_417/Y vdd NAND2X1
XAND2X2_28 AOI22X1_9/C INVX1_39/A gnd NOR2X1_27/B vdd AND2X2
XOAI21X1_267 INVX1_291/Y AOI22X1_86/Y AOI22X1_87/Y gnd OAI21X1_267/Y vdd OAI21X1
XNAND2X1_381 BUFX2_112/Y INVX1_433/Y gnd NAND2X1_381/Y vdd NAND2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_67/B gnd BUFX2_107/A vdd NOR2X1
XOAI21X1_231 INVX1_251/A INVX1_253/Y INVX1_252/Y gnd OAI21X1_231/Y vdd OAI21X1
XNAND2X1_345 INVX1_385/A BUFX2_38/Y gnd NAND2X1_345/Y vdd NAND2X1
XNOR2X1_31 gnd INVX1_47/Y gnd NOR2X1_31/Y vdd NOR2X1
XNAND3X1_177 NOR2X1_233/Y NAND3X1_176/Y OAI21X1_522/Y gnd NAND3X1_177/Y vdd NAND3X1
XINVX1_593 INVX1_96/A gnd INVX1_593/Y vdd INVX1
XOAI21X1_195 BUFX2_92/Y INVX1_209/Y OAI21X1_195/C gnd NAND3X1_69/C vdd OAI21X1
XNAND2X1_309 BUFX2_73/Y INVX1_345/A gnd OAI21X1_314/B vdd NAND2X1
XNOR2X1_228 NOR2X1_227/Y AND2X2_132/Y gnd INVX1_612/A vdd NOR2X1
XNAND3X1_141 NOR2X1_179/Y NAND3X1_140/Y NAND3X1_141/C gnd NAND3X1_141/Y vdd NAND3X1
XBUFX2_142 BUFX2_142/A gnd response_get[5] vdd BUFX2
XINVX1_557 INVX1_557/A gnd INVX1_557/Y vdd INVX1
XCLKBUF1_19 BUFX2_3/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XOAI21X1_159 INVX1_167/Y INVX1_170/Y AOI22X1_53/C gnd OAI21X1_159/Y vdd OAI21X1
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_192 NOR2X1_191/Y AND2X2_114/Y gnd INVX1_528/A vdd NOR2X1
XNAND2X1_273 INVX1_296/A NAND2X1_273/B gnd AOI22X1_89/A vdd NAND2X1
XBUFX2_106 BUFX2_103/A gnd INVX1_113/A vdd BUFX2
XINVX1_521 INVX1_437/A gnd INVX1_521/Y vdd INVX1
XDFFPOSX1_339 INVX1_578/A CLKBUF1_46/Y OAI21X1_514/Y gnd vdd DFFPOSX1
XNAND3X1_105 NOR2X1_125/Y NAND3X1_104/Y OAI21X1_306/Y gnd NAND3X1_105/Y vdd NAND3X1
XXNOR2X1_66 INVX1_237/A BUFX2_133/Y gnd XNOR2X1_66/Y vdd XNOR2X1
XOAI21X1_123 INVX1_129/Y NAND2X1_133/Y OAI21X1_123/C gnd DFFPOSX1_82/D vdd OAI21X1
XNOR2X1_156 NOR2X1_156/A AND2X2_96/Y gnd INVX1_444/A vdd NOR2X1
XNAND2X1_237 INVX1_251/A INVX1_254/Y gnd AOI22X1_76/D vdd NAND2X1
XDFFPOSX1_303 INVX1_515/A CLKBUF1_21/Y OAI21X1_460/Y gnd vdd DFFPOSX1
XINVX1_485 INVX1_485/A gnd INVX1_485/Y vdd INVX1
XXNOR2X1_30 BUFX2_17/Y INVX1_237/A gnd XNOR2X1_30/Y vdd XNOR2X1
XNOR2X1_120 NOR2X1_119/Y AND2X2_78/Y gnd AND2X2_84/B vdd NOR2X1
XNAND2X1_201 INVX1_209/A NAND2X1_9/B gnd NAND2X1_201/Y vdd NAND2X1
XFILL_4_1 gnd vdd FILL
XDFFPOSX1_267 INVX1_199/A CLKBUF1_6/Y OAI21X1_406/Y gnd vdd DFFPOSX1
XINVX1_449 AND2X2_8/Y gnd INVX1_449/Y vdd INVX1
XNAND2X1_165 INVX1_198/A INVX1_191/A gnd NOR2X1_67/A vdd NAND2X1
XDFFPOSX1_231 AND2X2_87/B CLKBUF1_41/Y OAI21X1_352/Y gnd vdd DFFPOSX1
XFILL_26_2 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XINVX1_413 INVX1_413/A gnd INVX1_413/Y vdd INVX1
XAOI21X1_63 INVX1_436/Y XNOR2X1_58/Y AOI21X1_63/C gnd AOI21X1_63/Y vdd AOI21X1
XFILL_16_2_1 gnd vdd FILL
XBUFX2_66 BUFX2_65/A gnd BUFX2_66/Y vdd BUFX2
XNAND2X1_129 NOR2X1_53/A BUFX2_105/Y gnd NAND2X1_129/Y vdd NAND2X1
XAOI21X1_27 INVX1_184/Y AOI21X1_27/B AOI21X1_27/C gnd AOI21X1_27/Y vdd AOI21X1
XINVX1_377 BUFX2_73/Y gnd INVX1_377/Y vdd INVX1
XDFFPOSX1_7 INVX1_22/A CLKBUF1_34/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XDFFPOSX1_195 INVX1_326/A CLKBUF1_3/Y OAI21X1_298/Y gnd vdd DFFPOSX1
XOAI21X1_556 INVX1_627/Y OAI21X1_556/B AOI22X1_183/Y gnd OAI21X1_556/Y vdd OAI21X1
XFILL_4_0_2 gnd vdd FILL
XBUFX2_30 RST_N gnd BUFX2_30/Y vdd BUFX2
XDFFPOSX1_93 INVX1_140/A CLKBUF1_8/Y NAND3X1_49/Y gnd vdd DFFPOSX1
XNAND2X1_90 INVX1_70/A BUFX2_43/Y gnd NAND2X1_90/Y vdd NAND2X1
XOAI21X1_75 INVX1_70/Y OAI21X1_75/B NOR2X1_37/Y gnd OAI21X1_75/Y vdd OAI21X1
XAOI22X1_161 AOI22X1_161/A AND2X2_126/Y AOI22X1_161/C NOR2X1_216/Y gnd AOI22X1_161/Y
+ vdd AOI22X1
XDFFPOSX1_159 AND2X2_65/B CLKBUF1_29/Y OAI21X1_242/Y gnd vdd DFFPOSX1
XOAI21X1_520 INVX1_585/Y AOI22X1_170/Y AOI22X1_171/Y gnd OAI21X1_520/Y vdd OAI21X1
XINVX1_341 INVX1_96/A gnd INVX1_341/Y vdd INVX1
XBUFX2_8 BUFX2_8/A gnd BUFX2_8/Y vdd BUFX2
XAOI22X1_68 INVX1_224/A INVX1_223/Y INVX1_225/Y AOI22X1_68/D gnd AOI22X1_68/Y vdd
+ AOI22X1
XNAND2X1_54 NAND2X1_54/A AOI22X1_9/Y gnd NAND2X1_54/Y vdd NAND2X1
XDFFPOSX1_123 INVX1_200/A CLKBUF1_49/Y OAI21X1_187/Y gnd vdd DFFPOSX1
XOAI21X1_39 NOR2X1_22/Y AOI21X1_4/Y BUFX2_139/A gnd NAND2X1_55/A vdd OAI21X1
XDFFPOSX1_57 INVX1_77/A CLKBUF1_51/Y NAND3X1_31/Y gnd vdd DFFPOSX1
XAOI22X1_125 AOI22X1_125/A AND2X2_99/Y OAI21X1_379/C NOR2X1_162/Y gnd OAI21X1_382/C
+ vdd AOI22X1
XOAI21X1_484 INVX1_543/Y OAI21X1_484/B OAI21X1_484/C gnd OAI21X1_484/Y vdd OAI21X1
XINVX1_305 AND2X2_72/B gnd INVX1_305/Y vdd INVX1
XAOI22X1_32 INVX1_98/A INVX1_97/Y INVX1_99/Y AOI22X1_32/D gnd AOI22X1_32/Y vdd AOI22X1
XFILL_25_0_0 gnd vdd FILL
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd BUFX2_22/A vdd NOR2X1
XFILL_3_3_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_23_2_1 gnd vdd FILL
XNAND2X1_18 INVX1_100/A INVX1_58/A gnd INVX1_7/A vdd NAND2X1
XDFFPOSX1_21 INVX1_32/A CLKBUF1_28/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XOAI21X1_448 INVX1_501/Y AOI22X1_146/Y OAI21X1_448/C gnd OAI21X1_448/Y vdd OAI21X1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XNAND3X1_95 NAND3X1_95/A NAND3X1_94/Y NAND3X1_95/C gnd NAND3X1_95/Y vdd NAND3X1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XOAI21X1_412 INVX1_459/Y AOI22X1_134/Y AOI22X1_135/Y gnd OAI21X1_412/Y vdd OAI21X1
XNAND2X1_526 AND2X2_20/A NAND2X1_526/B gnd NAND2X1_526/Y vdd NAND2X1
XNAND3X1_59 NOR2X1_70/Y NAND3X1_58/Y NAND3X1_59/C gnd NAND3X1_59/Y vdd NAND3X1
XNAND2X1_7 NAND2X1_7/A INVX1_170/A gnd NOR2X1_4/A vdd NAND2X1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd NOR2X1_77/B vdd INVX1
XOAI21X1_376 INVX1_417/Y OAI21X1_376/B OAI21X1_376/C gnd OAI21X1_376/Y vdd OAI21X1
XAND2X2_128 BUFX2_99/Y INVX1_479/A gnd AND2X2_128/Y vdd AND2X2
XNAND3X1_23 NOR2X1_31/Y NAND3X1_22/Y OAI21X1_53/Y gnd NAND3X1_23/Y vdd NAND3X1
XNAND2X1_490 INVX1_575/A INVX1_573/Y gnd OAI21X1_513/B vdd NAND2X1
XOAI21X1_340 INVX1_375/Y AOI22X1_110/Y OAI21X1_340/C gnd OAI21X1_340/Y vdd OAI21X1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XNAND2X1_454 INVX1_525/A INVX1_69/A gnd NAND2X1_454/Y vdd NAND2X1
XAND2X2_65 INVX1_251/A AND2X2_65/B gnd AND2X2_65/Y vdd AND2X2
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XOAI21X1_304 INVX1_333/Y AOI22X1_98/Y AOI22X1_99/Y gnd OAI21X1_304/Y vdd OAI21X1
XNAND2X1_418 BUFX2_134/Y INVX1_485/A gnd NAND2X1_418/Y vdd NAND2X1
XAND2X2_29 INVX1_42/A INVX1_51/A gnd INVX1_41/A vdd AND2X2
XNAND2X1_382 BUFX2_96/Y INVX1_436/Y gnd NAND2X1_382/Y vdd NAND2X1
XOAI21X1_268 INVX1_293/A INVX1_295/Y INVX1_294/Y gnd OAI21X1_268/Y vdd OAI21X1
XFILL_17_1 gnd vdd FILL
XNOR2X1_68 gnd INVX1_166/Y gnd NOR2X1_68/Y vdd NOR2X1
XOAI21X1_232 BUFX2_95/Y INVX1_251/Y OAI21X1_231/Y gnd NAND3X1_81/C vdd OAI21X1
XNAND2X1_346 INVX1_387/A NAND2X1_345/Y gnd AOI22X1_115/A vdd NAND2X1
XNAND3X1_178 BUFX2_78/Y INVX1_596/Y INVX1_597/Y gnd NAND3X1_179/B vdd NAND3X1
XNOR2X1_32 INVX1_4/A INVX1_50/Y gnd NOR2X1_32/Y vdd NOR2X1
XINVX1_594 BUFX2_78/Y gnd INVX1_594/Y vdd INVX1
XOAI21X1_196 INVX1_209/Y INVX1_212/Y AOI22X1_65/C gnd OAI21X1_197/C vdd OAI21X1
XNOR2X1_229 INVX1_606/A INVX1_592/A gnd NOR2X1_229/Y vdd NOR2X1
XNAND2X1_310 AND2X2_85/A INVX1_342/Y gnd OAI21X1_315/B vdd NAND2X1
XINVX1_558 BUFX2_34/Y gnd INVX1_558/Y vdd INVX1
XBUFX2_143 BUFX2_143/A gnd response_get[6] vdd BUFX2
XCLKBUF1_20 BUFX2_6/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XNAND3X1_142 BUFX2_90/Y INVX1_470/Y INVX1_471/Y gnd NAND3X1_142/Y vdd NAND3X1
XOAI21X1_160 INVX1_171/Y NAND2X1_167/Y OAI21X1_159/Y gnd OAI21X1_160/Y vdd OAI21X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_193 INVX1_522/A INVX1_508/A gnd NOR2X1_193/Y vdd NOR2X1
XNAND2X1_274 BUFX2_51/Y AND2X2_71/B gnd NAND2X1_274/Y vdd NAND2X1
XDFFPOSX1_340 INVX1_576/A CLKBUF1_38/Y AOI21X1_83/Y gnd vdd DFFPOSX1
XBUFX2_107 BUFX2_107/A gnd INVX1_204/A vdd BUFX2
XNAND3X1_106 BUFX2_77/Y INVX1_344/Y INVX1_345/Y gnd NAND3X1_106/Y vdd NAND3X1
XINVX1_522 INVX1_522/A gnd INVX1_522/Y vdd INVX1
XXNOR2X1_67 INVX1_498/A BUFX2_130/Y gnd AOI21X1_72/B vdd XNOR2X1
XOAI21X1_124 INVX1_126/Y NAND2X1_134/Y NOR2X1_55/Y gnd AOI21X1_19/C vdd OAI21X1
XNOR2X1_157 AND2X2_96/A AND2X2_98/B gnd NOR2X1_157/Y vdd NOR2X1
XNAND2X1_238 NOR2X1_95/A BUFX2_95/Y gnd NAND2X1_239/B vdd NAND2X1
XINVX1_486 INVX1_486/A gnd INVX1_486/Y vdd INVX1
XDFFPOSX1_304 INVX1_513/A CLKBUF1_21/Y AOI21X1_74/Y gnd vdd DFFPOSX1
XXNOR2X1_31 BUFX2_15/Y INVX1_244/A gnd XNOR2X1_31/Y vdd XNOR2X1
XNOR2X1_121 INVX1_354/A AND2X2_79/B gnd NOR2X1_122/A vdd NOR2X1
XFILL_10_3_0 gnd vdd FILL
XNAND2X1_202 BUFX2_92/Y INVX1_209/Y gnd OAI21X1_198/B vdd NAND2X1
XDFFPOSX1_268 AND2X2_8/A CLKBUF1_6/Y AOI21X1_65/Y gnd vdd DFFPOSX1
XINVX1_450 AND2X2_8/A gnd INVX1_450/Y vdd INVX1
XNAND2X1_166 NOR2X1_73/A INVX1_205/A gnd NOR2X1_67/B vdd NAND2X1
XAOI21X1_64 INVX1_443/Y AOI21X1_64/B AOI21X1_64/C gnd AOI21X1_64/Y vdd AOI21X1
XDFFPOSX1_232 INVX1_387/A CLKBUF1_41/Y AOI21X1_56/Y gnd vdd DFFPOSX1
XFILL_18_0_1 gnd vdd FILL
XINVX1_414 AND2X2_6/Y gnd INVX1_414/Y vdd INVX1
XFILL_16_2_2 gnd vdd FILL
XBUFX2_67 BUFX2_67/A gnd BUFX2_67/Y vdd BUFX2
XNAND2X1_130 INVX1_121/A NAND2X1_129/Y gnd AOI22X1_39/A vdd NAND2X1
XAOI21X1_28 INVX1_191/Y XNOR2X1_23/Y AOI21X1_28/C gnd AOI21X1_28/Y vdd AOI21X1
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XDFFPOSX1_8 INVX1_23/A CLKBUF1_18/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_196 INVX1_324/A CLKBUF1_40/Y AOI21X1_47/Y gnd vdd DFFPOSX1
XBUFX2_31 RST_N gnd BUFX2_31/Y vdd BUFX2
XDFFPOSX1_94 AOI22X1_47/C CLKBUF1_43/Y OAI21X1_142/Y gnd vdd DFFPOSX1
XDFFPOSX1_160 AND2X2_64/B CLKBUF1_37/Y AOI21X1_38/Y gnd vdd DFFPOSX1
XNAND2X1_91 INVX1_72/A NAND2X1_90/Y gnd NAND2X1_91/Y vdd NAND2X1
XOAI21X1_76 INVX1_74/Y OAI21X1_76/B OAI21X1_76/C gnd OAI21X1_76/Y vdd OAI21X1
XAOI22X1_162 INVX1_553/A INVX1_552/Y INVX1_554/Y NAND2X1_476/Y gnd OAI21X1_496/B vdd
+ AOI22X1
XINVX1_342 BUFX2_77/Y gnd INVX1_342/Y vdd INVX1
XOAI21X1_521 BUFX2_24/Y INVX1_589/Y INVX1_588/Y gnd OAI21X1_521/Y vdd OAI21X1
XBUFX2_9 BUFX2_8/A gnd BUFX2_9/Y vdd BUFX2
XFILL_17_3_0 gnd vdd FILL
XAOI22X1_69 AOI22X1_69/A AND2X2_60/Y AOI22X1_69/C NOR2X1_86/Y gnd AOI22X1_69/Y vdd
+ AOI22X1
XNAND2X1_55 NAND2X1_55/A AOI22X1_10/Y gnd NAND2X1_55/Y vdd NAND2X1
XDFFPOSX1_124 INVX1_198/A CLKBUF1_49/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XAOI22X1_126 INVX1_427/A INVX1_426/Y INVX1_428/Y NAND2X1_377/Y gnd AOI22X1_126/Y vdd
+ AOI22X1
XOAI21X1_40 NOR2X1_22/Y AOI21X1_4/Y BUFX2_140/A gnd NAND2X1_56/A vdd OAI21X1
XDFFPOSX1_58 OAI21X1_85/C CLKBUF1_3/Y OAI21X1_86/Y gnd vdd DFFPOSX1
XINVX1_306 INVX1_96/A gnd INVX1_306/Y vdd INVX1
XOAI21X1_485 BUFX2_74/Y INVX1_547/Y INVX1_546/Y gnd OAI21X1_486/C vdd OAI21X1
XAOI22X1_33 AOI22X1_33/A AND2X2_39/Y AOI22X1_33/C NOR2X1_47/Y gnd AOI22X1_33/Y vdd
+ AOI22X1
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd BUFX2_73/A vdd NOR2X1
XFILL_25_0_1 gnd vdd FILL
XFILL_23_2_2 gnd vdd FILL
XFILL_3_3_2 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XDFFPOSX1_22 INVX1_33/A CLKBUF1_13/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XNAND2X1_19 INVX1_268/A INVX1_226/A gnd NOR2X1_9/B vdd NAND2X1
XOAI21X1_449 BUFX2_25/Y INVX1_505/Y INVX1_504/Y gnd OAI21X1_449/Y vdd OAI21X1
XINVX1_270 INVX1_39/A gnd INVX1_270/Y vdd INVX1
XNAND3X1_96 BUFX2_18/Y INVX1_309/Y INVX1_310/Y gnd NAND3X1_97/B vdd NAND3X1
XINVX1_234 INVX1_417/A gnd INVX1_234/Y vdd INVX1
XOAI21X1_413 BUFX2_83/Y INVX1_463/Y INVX1_462/Y gnd OAI21X1_414/C vdd OAI21X1
XNAND3X1_60 BUFX2_108/Y NOR2X1_73/B INVX1_184/Y gnd NAND3X1_60/Y vdd NAND3X1
XNAND2X1_527 BUFX2_10/Y AND2X2_21/A gnd NAND2X1_527/Y vdd NAND2X1
XNAND2X1_8 NAND2X1_8/A INVX1_427/A gnd NOR2X1_4/B vdd NAND2X1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XOAI21X1_377 BUFX2_80/Y INVX1_421/Y INVX1_420/Y gnd OAI21X1_377/Y vdd OAI21X1
XFILL_24_3_0 gnd vdd FILL
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XAND2X2_129 INVX1_547/A INVX1_570/A gnd AND2X2_129/Y vdd AND2X2
XNAND3X1_24 INVX1_55/A INVX1_57/Y INVX1_58/Y gnd NAND3X1_25/B vdd NAND3X1
XNAND2X1_491 BUFX2_124/Y INVX1_576/Y gnd NAND2X1_491/Y vdd NAND2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_162 BUFX2_48/Y gnd INVX1_162/Y vdd INVX1
XOAI21X1_341 BUFX2_75/Y INVX1_379/Y INVX1_378/Y gnd OAI21X1_342/C vdd OAI21X1
XNAND2X1_455 AND2X2_13/A NAND2X1_454/Y gnd NAND2X1_455/Y vdd NAND2X1
XAND2X2_66 BUFX2_51/Y AND2X2_66/B gnd AND2X2_66/Y vdd AND2X2
XOAI21X1_305 BUFX2_22/Y INVX1_337/Y INVX1_336/Y gnd OAI21X1_306/C vdd OAI21X1
XINVX1_126 NOR2X1_56/A gnd INVX1_126/Y vdd INVX1
XNAND2X1_419 INVX1_484/A INVX1_482/Y gnd OAI21X1_435/B vdd NAND2X1
XAND2X2_30 INVX1_41/A INVX1_45/A gnd AND2X2_30/Y vdd AND2X2
XOAI21X1_269 BUFX2_100/Y INVX1_293/Y OAI21X1_268/Y gnd NAND3X1_93/C vdd OAI21X1
XNAND2X1_383 INVX1_434/A INVX1_421/A gnd NAND2X1_383/Y vdd NAND2X1
XNOR2X1_69 INVX1_168/A INVX1_169/Y gnd NOR2X1_69/Y vdd NOR2X1
XOAI21X1_233 INVX1_251/Y INVX1_254/Y AOI22X1_77/C gnd OAI21X1_234/C vdd OAI21X1
XNAND2X1_347 BUFX2_88/Y INVX1_394/A gnd NAND2X1_347/Y vdd NAND2X1
XNAND3X1_179 NOR2X1_235/Y NAND3X1_179/B NAND3X1_179/C gnd NAND3X1_179/Y vdd NAND3X1
XINVX1_595 NAND2X1_6/B gnd INVX1_595/Y vdd INVX1
XNOR2X1_33 gnd INVX1_54/Y gnd NOR2X1_33/Y vdd NOR2X1
XNAND2X1_311 BUFX2_77/Y INVX1_345/Y gnd NAND2X1_311/Y vdd NAND2X1
XOAI21X1_197 INVX1_213/Y NAND2X1_201/Y OAI21X1_197/C gnd OAI21X1_197/Y vdd OAI21X1
XNOR2X1_230 NOR2X1_229/Y NOR2X1_230/B gnd INVX1_619/A vdd NOR2X1
XINVX1_559 BUFX2_98/Y gnd INVX1_559/Y vdd INVX1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XCLKBUF1_21 BUFX2_4/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XNAND3X1_143 NOR2X1_181/Y NAND3X1_142/Y OAI21X1_420/Y gnd NAND3X1_143/Y vdd NAND3X1
XOAI21X1_161 INVX1_168/Y NAND2X1_168/Y NOR2X1_68/Y gnd AOI21X1_25/C vdd OAI21X1
XFILL_11_0_2 gnd vdd FILL
XNOR2X1_194 NOR2X1_193/Y AND2X2_115/Y gnd INVX1_535/A vdd NOR2X1
XNAND2X1_275 INVX1_293/A INVX1_300/Y gnd NAND2X1_275/Y vdd NAND2X1
XDFFPOSX1_341 INVX1_574/A CLKBUF1_38/Y NAND3X1_173/Y gnd vdd DFFPOSX1
XBUFX2_108 BUFX2_107/A gnd BUFX2_108/Y vdd BUFX2
XINVX1_523 BUFX2_32/Y gnd INVX1_523/Y vdd INVX1
XNAND3X1_107 NOR2X1_127/Y NAND3X1_106/Y NAND3X1_107/C gnd NAND3X1_107/Y vdd NAND3X1
XNOR2X1_158 NOR2X1_157/Y AND2X2_97/Y gnd INVX1_451/A vdd NOR2X1
XOAI21X1_125 INVX1_130/Y AOI22X1_40/Y AOI22X1_41/Y gnd OAI21X1_125/Y vdd OAI21X1
XXNOR2X1_68 BUFX2_61/Y INVX1_43/A gnd XNOR2X1_68/Y vdd XNOR2X1
XNAND2X1_239 INVX1_254/A NAND2X1_239/B gnd AOI22X1_77/A vdd NAND2X1
XINVX1_487 INVX1_487/A gnd INVX1_487/Y vdd INVX1
XDFFPOSX1_305 INVX1_511/A CLKBUF1_21/Y NAND3X1_155/Y gnd vdd DFFPOSX1
XXNOR2X1_32 BUFX2_95/Y INVX1_251/A gnd AOI21X1_37/B vdd XNOR2X1
XNOR2X1_122 NOR2X1_122/A AND2X2_79/Y gnd INVX1_367/A vdd NOR2X1
XNAND2X1_203 INVX1_209/A INVX1_212/Y gnd AOI22X1_64/D vdd NAND2X1
XDFFPOSX1_269 INVX1_448/A CLKBUF1_6/Y NAND3X1_137/Y gnd vdd DFFPOSX1
XFILL_10_3_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XINVX1_451 INVX1_451/A gnd INVX1_451/Y vdd INVX1
XNAND2X1_167 INVX1_167/A INVX1_170/A gnd NAND2X1_167/Y vdd NAND2X1
XAOI21X1_65 INVX1_450/Y AOI21X1_65/B AOI21X1_65/C gnd AOI21X1_65/Y vdd AOI21X1
XINVX1_415 AND2X2_6/A gnd INVX1_415/Y vdd INVX1
XDFFPOSX1_233 INVX1_385/A CLKBUF1_41/Y NAND3X1_119/Y gnd vdd DFFPOSX1
XFILL_18_0_2 gnd vdd FILL
XBUFX2_68 BUFX2_67/A gnd BUFX2_68/Y vdd BUFX2
XNAND2X1_131 INVX1_156/A INVX1_149/A gnd NOR2X1_54/A vdd NAND2X1
XDFFPOSX1_9 INVX1_24/A CLKBUF1_18/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XAOI21X1_29 INVX1_198/Y AOI21X1_29/B AOI21X1_29/C gnd AOI21X1_29/Y vdd AOI21X1
XINVX1_379 BUFX2_37/Y gnd INVX1_379/Y vdd INVX1
XDFFPOSX1_197 AND2X2_18/B CLKBUF1_44/Y NAND3X1_101/Y gnd vdd DFFPOSX1
XBUFX2_32 RST_N gnd BUFX2_32/Y vdd BUFX2
XNAND2X1_92 INVX1_76/A INVX1_79/A gnd OAI21X1_80/B vdd NAND2X1
XDFFPOSX1_95 INVX1_151/A CLKBUF1_43/Y OAI21X1_144/Y gnd vdd DFFPOSX1
XOAI21X1_77 INVX1_76/A INVX1_78/Y INVX1_77/Y gnd OAI21X1_77/Y vdd OAI21X1
XDFFPOSX1_161 NOR2X1_97/A CLKBUF1_29/Y NAND3X1_83/Y gnd vdd DFFPOSX1
XAOI22X1_163 AOI22X1_163/A AND2X2_127/Y OAI21X1_493/C NOR2X1_218/Y gnd OAI21X1_496/C
+ vdd AOI22X1
XINVX1_343 INVX1_343/A gnd INVX1_343/Y vdd INVX1
XOAI21X1_522 BUFX2_12/Y INVX1_587/Y OAI21X1_521/Y gnd OAI21X1_522/Y vdd OAI21X1
XFILL_19_1_0 gnd vdd FILL
XAOI22X1_70 AND2X2_6/B INVX1_230/Y NOR2X1_88/B AOI22X1_70/D gnd AOI22X1_70/Y vdd AOI22X1
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_41 NOR2X1_22/Y AOI21X1_4/Y BUFX2_141/A gnd NAND2X1_57/A vdd OAI21X1
XNAND2X1_56 NAND2X1_56/A AOI22X1_11/Y gnd NAND2X1_56/Y vdd NAND2X1
XDFFPOSX1_125 AND2X2_8/B CLKBUF1_6/Y NAND3X1_65/Y gnd vdd DFFPOSX1
XAOI22X1_127 NAND2X1_379/Y AND2X2_100/Y OAI21X1_385/C NOR2X1_164/Y gnd AOI22X1_127/Y
+ vdd AOI22X1
XINVX1_307 BUFX2_18/Y gnd INVX1_307/Y vdd INVX1
XDFFPOSX1_59 INVX1_88/A CLKBUF1_48/Y OAI21X1_88/Y gnd vdd DFFPOSX1
XOAI21X1_486 INVX1_547/A INVX1_545/Y OAI21X1_486/C gnd NAND3X1_165/C vdd OAI21X1
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd BUFX2_79/A vdd NOR2X1
XAOI22X1_34 AND2X2_2/B INVX1_104/Y NOR2X1_49/B AOI22X1_34/D gnd AOI22X1_34/Y vdd AOI22X1
XFILL_25_0_2 gnd vdd FILL
XFILL_5_1_2 gnd vdd FILL
XDFFPOSX1_23 INVX1_34/A CLKBUF1_20/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XNAND2X1_20 INVX1_28/A INVX1_310/A gnd NOR2X1_11/A vdd NAND2X1
XINVX1_271 BUFX2_33/Y gnd INVX1_271/Y vdd INVX1
XOAI21X1_450 BUFX2_61/Y INVX1_503/Y OAI21X1_449/Y gnd NAND3X1_153/C vdd OAI21X1
XNAND3X1_97 NOR2X1_111/Y NAND3X1_97/B NAND3X1_97/C gnd NAND3X1_97/Y vdd NAND3X1
XNAND3X1_61 NOR2X1_72/Y NAND3X1_60/Y NAND3X1_61/C gnd NAND3X1_61/Y vdd NAND3X1
XINVX1_235 INVX1_235/A gnd INVX1_235/Y vdd INVX1
XOAI21X1_414 INVX1_463/A INVX1_461/Y OAI21X1_414/C gnd NAND3X1_141/C vdd OAI21X1
XNAND2X1_9 INVX1_392/A NAND2X1_9/B gnd NOR2X1_5/A vdd NAND2X1
XNAND2X1_528 INVX1_624/A INVX1_622/Y gnd NAND2X1_528/Y vdd NAND2X1
XFILL_26_1_0 gnd vdd FILL
XFILL_24_3_1 gnd vdd FILL
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XFILL_6_2_0 gnd vdd FILL
XOAI21X1_378 INVX1_421/A INVX1_419/Y OAI21X1_377/Y gnd OAI21X1_378/Y vdd OAI21X1
XAND2X2_130 INVX1_554/A INVX1_577/A gnd AND2X2_130/Y vdd AND2X2
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XNAND3X1_25 NOR2X1_33/Y NAND3X1_25/B NAND3X1_25/C gnd NAND3X1_25/Y vdd NAND3X1
XNAND2X1_492 INVX1_574/A INVX1_575/A gnd NAND2X1_493/B vdd NAND2X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XOAI21X1_342 BUFX2_38/Y INVX1_377/Y OAI21X1_342/C gnd OAI21X1_342/Y vdd OAI21X1
XNAND2X1_456 BUFX2_62/Y AND2X2_14/A gnd NAND2X1_456/Y vdd NAND2X1
XAND2X2_67 BUFX2_58/Y INVX1_269/A gnd AND2X2_67/Y vdd AND2X2
XINVX1_127 BUFX2_82/Y gnd NOR2X1_56/B vdd INVX1
XNAND2X1_420 BUFX2_134/Y INVX1_485/Y gnd NAND2X1_420/Y vdd NAND2X1
XOAI21X1_306 BUFX2_117/Y INVX1_335/Y OAI21X1_306/C gnd OAI21X1_306/Y vdd OAI21X1
XAND2X2_31 BUFX2_56/Y INVX1_52/A gnd AND2X2_31/Y vdd AND2X2
XOAI21X1_270 INVX1_293/Y INVX1_296/Y AOI22X1_89/C gnd OAI21X1_271/C vdd OAI21X1
XNAND2X1_384 INVX1_436/A NAND2X1_383/Y gnd NAND2X1_384/Y vdd NAND2X1
XNOR2X1_70 gnd NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XOAI21X1_234 INVX1_255/Y NAND2X1_235/Y OAI21X1_234/C gnd OAI21X1_234/Y vdd OAI21X1
XNAND2X1_348 BUFX2_36/Y INVX1_391/Y gnd OAI21X1_357/B vdd NAND2X1
XNAND3X1_180 BUFX2_99/Y INVX1_603/Y INVX1_604/Y gnd NAND3X1_181/B vdd NAND3X1
XINVX1_596 BUFX2_13/Y gnd INVX1_596/Y vdd INVX1
XOAI21X1_198 INVX1_210/Y OAI21X1_198/B NOR2X1_81/Y gnd AOI21X1_31/C vdd OAI21X1
XNOR2X1_34 INVX1_56/A INVX1_57/Y gnd NOR2X1_34/Y vdd NOR2X1
XNAND2X1_312 INVX1_343/A AND2X2_85/A gnd NAND2X1_313/B vdd NAND2X1
XNOR2X1_231 INVX1_599/A INVX1_592/A gnd NOR2X1_232/A vdd NOR2X1
XNAND3X1_144 BUFX2_98/Y INVX1_477/Y INVX1_478/Y gnd NAND3X1_144/Y vdd NAND3X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX1_560 INVX1_560/A gnd INVX1_560/Y vdd INVX1
XCLKBUF1_22 BUFX2_4/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XOAI21X1_162 INVX1_172/Y AOI22X1_52/Y AOI22X1_53/Y gnd OAI21X1_162/Y vdd OAI21X1
XNOR2X1_195 INVX1_515/A INVX1_508/A gnd NOR2X1_195/Y vdd NOR2X1
XNAND2X1_276 BUFX2_52/Y INVX1_303/Y gnd AOI22X1_90/D vdd NAND2X1
XBUFX2_109 BUFX2_107/A gnd INVX1_197/A vdd BUFX2
XNAND3X1_108 BUFX2_86/Y INVX1_351/Y INVX1_352/Y gnd NAND3X1_109/B vdd NAND3X1
XINVX1_524 BUFX2_66/Y gnd INVX1_524/Y vdd INVX1
XDFFPOSX1_342 OAI21X1_517/C CLKBUF1_9/Y OAI21X1_518/Y gnd vdd DFFPOSX1
XXNOR2X1_69 BUFX2_63/Y BUFX2_89/Y gnd XNOR2X1_69/Y vdd XNOR2X1
XNOR2X1_159 INVX1_431/A AND2X2_98/B gnd NOR2X1_159/Y vdd NOR2X1
XOAI21X1_126 BUFX2_50/Y NOR2X1_58/B INVX1_133/Y gnd OAI21X1_126/Y vdd OAI21X1
XNAND2X1_240 BUFX2_52/Y AND2X2_64/B gnd NAND2X1_240/Y vdd NAND2X1
XINVX1_488 BUFX2_34/Y gnd INVX1_488/Y vdd INVX1
XDFFPOSX1_306 AOI22X1_153/C CLKBUF1_29/Y OAI21X1_464/Y gnd vdd DFFPOSX1
XXNOR2X1_33 INVX1_251/A BUFX2_52/Y gnd AOI21X1_38/B vdd XNOR2X1
XFILL_12_1_1 gnd vdd FILL
XNOR2X1_123 AND2X2_80/A AND2X2_79/B gnd NOR2X1_123/Y vdd NOR2X1
XNAND2X1_204 INVX1_210/A BUFX2_92/Y gnd NAND2X1_205/B vdd NAND2X1
XDFFPOSX1_270 OAI21X1_409/C CLKBUF1_45/Y OAI21X1_410/Y gnd vdd DFFPOSX1
XFILL_10_3_2 gnd vdd FILL
XINVX1_452 INVX1_199/A gnd INVX1_452/Y vdd INVX1
XNAND2X1_168 BUFX2_85/Y INVX1_167/Y gnd NAND2X1_168/Y vdd NAND2X1
XINVX1_416 INVX1_416/A gnd INVX1_416/Y vdd INVX1
XAOI21X1_66 INVX1_457/Y XNOR2X1_61/Y AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XDFFPOSX1_234 AOI22X1_117/C CLKBUF1_44/Y OAI21X1_356/Y gnd vdd DFFPOSX1
XBUFX2_69 BUFX2_67/A gnd BUFX2_69/Y vdd BUFX2
XNAND2X1_132 INVX1_140/A INVX1_163/A gnd NOR2X1_54/B vdd NAND2X1
XDFFPOSX1_198 AOI22X1_99/C CLKBUF1_7/Y OAI21X1_302/Y gnd vdd DFFPOSX1
XAOI21X1_30 INVX1_205/Y XNOR2X1_25/Y AOI21X1_30/C gnd AOI21X1_30/Y vdd AOI21X1
XINVX1_380 INVX1_380/A gnd INVX1_380/Y vdd INVX1
XBUFX2_33 RST_N gnd BUFX2_33/Y vdd BUFX2
XOAI21X1_78 BUFX2_42/Y INVX1_76/Y OAI21X1_77/Y gnd OAI21X1_78/Y vdd OAI21X1
XNAND2X1_93 BUFX2_42/Y INVX1_76/Y gnd OAI21X1_81/B vdd NAND2X1
XDFFPOSX1_96 INVX1_149/A CLKBUF1_27/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XAOI22X1_164 INVX1_560/A INVX1_559/Y INVX1_561/Y AOI22X1_164/D gnd OAI21X1_502/B vdd
+ AOI22X1
XINVX1_344 AND2X2_85/A gnd INVX1_344/Y vdd INVX1
XDFFPOSX1_162 AOI22X1_81/C CLKBUF1_46/Y OAI21X1_246/Y gnd vdd DFFPOSX1
XFILL_1_0_0 gnd vdd FILL
XOAI21X1_523 INVX1_587/Y INVX1_590/Y AOI22X1_173/C gnd OAI21X1_524/C vdd OAI21X1
XFILL_19_1_1 gnd vdd FILL
XAOI22X1_71 AOI22X1_71/A AND2X2_61/Y AOI22X1_71/C NOR2X1_88/Y gnd AOI22X1_71/Y vdd
+ AOI22X1
XFILL_17_3_2 gnd vdd FILL
XNAND2X1_57 NAND2X1_57/A NAND2X1_57/B gnd NAND2X1_57/Y vdd NAND2X1
XOAI21X1_42 NOR2X1_22/Y AOI21X1_4/Y BUFX2_142/A gnd NAND2X1_58/A vdd OAI21X1
XDFFPOSX1_60 INVX1_86/A CLKBUF1_48/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 AOI22X1_63/C CLKBUF1_16/Y OAI21X1_191/Y gnd vdd DFFPOSX1
XAOI22X1_128 INVX1_434/A INVX1_433/Y INVX1_435/Y NAND2X1_382/Y gnd OAI21X1_394/B vdd
+ AOI22X1
XOAI21X1_487 INVX1_545/Y INVX1_548/Y AOI22X1_161/C gnd OAI21X1_488/C vdd OAI21X1
XINVX1_308 INVX1_308/A gnd INVX1_308/Y vdd INVX1
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd BUFX2_85/A vdd NOR2X1
XAOI22X1_35 AOI22X1_35/A AND2X2_40/Y AOI22X1_35/C NOR2X1_49/Y gnd AOI22X1_35/Y vdd
+ AOI22X1
XNAND2X1_21 INVX1_184/A INVX1_142/A gnd NOR2X1_11/B vdd NAND2X1
XFILL_8_1 gnd vdd FILL
XDFFPOSX1_24 INVX1_35/A CLKBUF1_13/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XINVX1_272 AND2X2_9/Y gnd INVX1_272/Y vdd INVX1
XOAI21X1_451 INVX1_503/Y INVX1_506/Y AOI22X1_149/C gnd OAI21X1_451/Y vdd OAI21X1
XNAND3X1_98 INVX1_498/A INVX1_316/Y INVX1_317/Y gnd NAND3X1_98/Y vdd NAND3X1
XINVX1_236 BUFX2_34/Y gnd INVX1_236/Y vdd INVX1
XOAI21X1_415 INVX1_461/Y INVX1_464/Y AOI22X1_137/C gnd OAI21X1_416/C vdd OAI21X1
XNAND3X1_62 AND2X2_3/Y NOR2X1_75/B INVX1_191/Y gnd NAND3X1_62/Y vdd NAND3X1
XNAND2X1_529 BUFX2_10/Y INVX1_625/Y gnd AOI22X1_182/D vdd NAND2X1
XFILL_6_2_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XFILL_24_3_2 gnd vdd FILL
XINVX1_82 INVX1_96/A gnd INVX1_82/Y vdd INVX1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XOAI21X1_379 INVX1_419/Y INVX1_422/Y OAI21X1_379/C gnd OAI21X1_380/C vdd OAI21X1
XAND2X2_131 INVX1_580/A INVX1_584/A gnd AND2X2_131/Y vdd AND2X2
XNAND3X1_26 AND2X2_1/Y INVX1_64/Y INVX1_65/Y gnd NAND3X1_26/Y vdd NAND3X1
XNAND2X1_493 INVX1_576/A NAND2X1_493/B gnd AOI22X1_169/A vdd NAND2X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_164 AND2X2_49/B gnd INVX1_164/Y vdd INVX1
XOAI21X1_343 INVX1_377/Y INVX1_380/Y AOI22X1_113/C gnd OAI21X1_343/Y vdd OAI21X1
XNAND2X1_457 INVX1_244/A INVX1_531/Y gnd OAI21X1_477/B vdd NAND2X1
XAND2X2_68 AND2X2_9/Y INVX1_459/A gnd AND2X2_68/Y vdd AND2X2
XINVX1_128 NAND2X1_5/B gnd INVX1_128/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XOAI21X1_307 INVX1_335/Y INVX1_338/Y OAI21X1_307/C gnd OAI21X1_308/C vdd OAI21X1
XNAND2X1_421 INVX1_483/A INVX1_484/A gnd NAND2X1_421/Y vdd NAND2X1
XAND2X2_32 BUFX2_43/Y INVX1_59/A gnd AND2X2_32/Y vdd AND2X2
XOAI21X1_271 INVX1_297/Y OAI21X1_271/B OAI21X1_271/C gnd OAI21X1_271/Y vdd OAI21X1
XNAND2X1_385 INVX1_440/A AND2X2_7/A gnd NAND2X1_385/Y vdd NAND2X1
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XOAI21X1_235 INVX1_252/Y NAND2X1_236/Y NOR2X1_94/Y gnd AOI21X1_37/C vdd OAI21X1
XNAND2X1_349 BUFX2_88/Y INVX1_394/Y gnd AOI22X1_116/D vdd NAND2X1
XNAND3X1_181 NOR2X1_237/Y NAND3X1_181/B NAND3X1_181/C gnd NAND3X1_181/Y vdd NAND3X1
XINVX1_597 INVX1_597/A gnd INVX1_597/Y vdd INVX1
XOAI21X1_199 INVX1_214/Y AOI22X1_64/Y AOI22X1_65/Y gnd OAI21X1_199/Y vdd OAI21X1
XNOR2X1_35 gnd INVX1_61/Y gnd NOR2X1_35/Y vdd NOR2X1
XNAND2X1_313 INVX1_345/A NAND2X1_313/B gnd AOI22X1_103/A vdd NAND2X1
XNOR2X1_232 NOR2X1_232/A AND2X2_134/Y gnd INVX1_626/A vdd NOR2X1
XNAND3X1_145 NOR2X1_183/Y NAND3X1_144/Y OAI21X1_426/Y gnd NAND3X1_145/Y vdd NAND3X1
XCLKBUF1_23 BUFX2_2/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XINVX1_561 BUFX2_125/Y gnd INVX1_561/Y vdd INVX1
XOR2X2_3 OR2X2_5/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XOAI21X1_163 BUFX2_54/Y NOR2X1_71/B INVX1_175/Y gnd OAI21X1_164/C vdd OAI21X1
XNOR2X1_196 NOR2X1_195/Y NOR2X1_196/B gnd INVX1_542/A vdd NOR2X1
XNAND2X1_277 INVX1_301/A INVX1_293/A gnd NAND2X1_277/Y vdd NAND2X1
XBUFX2_110 BUFX2_107/A gnd INVX1_190/A vdd BUFX2
XNAND3X1_109 NOR2X1_129/Y NAND3X1_109/B NAND3X1_109/C gnd NAND3X1_109/Y vdd NAND3X1
XINVX1_525 INVX1_525/A gnd INVX1_525/Y vdd INVX1
XDFFPOSX1_343 INVX1_325/A CLKBUF1_25/Y OAI21X1_520/Y gnd vdd DFFPOSX1
XOAI21X1_127 INVX1_125/A INVX1_132/Y OAI21X1_126/Y gnd NAND3X1_47/C vdd OAI21X1
XXNOR2X1_70 BUFX2_65/Y BUFX2_93/Y gnd XNOR2X1_70/Y vdd XNOR2X1
XNOR2X1_160 NOR2X1_159/Y AND2X2_98/Y gnd INVX1_458/A vdd NOR2X1
XNAND2X1_241 INVX1_251/A INVX1_258/Y gnd OAI21X1_241/B vdd NAND2X1
XDFFPOSX1_307 INVX1_522/A CLKBUF1_25/Y OAI21X1_466/Y gnd vdd DFFPOSX1
XINVX1_489 BUFX2_129/Y gnd INVX1_489/Y vdd INVX1
XFILL_21_1 gnd vdd FILL
XXNOR2X1_34 BUFX2_68/Y BUFX2_60/Y gnd AOI21X1_39/B vdd XNOR2X1
XFILL_12_1_2 gnd vdd FILL
XNOR2X1_124 NOR2X1_123/Y AND2X2_80/Y gnd AND2X2_86/B vdd NOR2X1
XNAND2X1_205 NAND2X1_9/B NAND2X1_205/B gnd AOI22X1_65/A vdd NAND2X1
XINVX1_453 BUFX2_31/Y gnd INVX1_453/Y vdd INVX1
XDFFPOSX1_271 INVX1_459/A CLKBUF1_13/Y OAI21X1_412/Y gnd vdd DFFPOSX1
XNAND2X1_169 INVX1_167/A INVX1_170/Y gnd AOI22X1_52/D vdd NAND2X1
XINVX1_417 INVX1_417/A gnd INVX1_417/Y vdd INVX1
XAOI21X1_67 INVX1_464/Y XNOR2X1_62/Y AOI21X1_67/C gnd AOI21X1_67/Y vdd AOI21X1
XDFFPOSX1_235 AND2X2_88/A CLKBUF1_7/Y OAI21X1_358/Y gnd vdd DFFPOSX1
XBUFX2_70 BUFX2_67/A gnd BUFX2_70/Y vdd BUFX2
XNAND2X1_133 INVX1_125/A NAND2X1_5/B gnd NAND2X1_133/Y vdd NAND2X1
XFILL_13_2_0 gnd vdd FILL
XAOI21X1_31 INVX1_212/Y XNOR2X1_26/Y AOI21X1_31/C gnd AOI21X1_31/Y vdd AOI21X1
XDFFPOSX1_199 INVX1_333/A CLKBUF1_3/Y OAI21X1_304/Y gnd vdd DFFPOSX1
XINVX1_381 INVX1_88/A gnd INVX1_381/Y vdd INVX1
XBUFX2_34 RST_N gnd BUFX2_34/Y vdd BUFX2
XDFFPOSX1_97 AND2X2_5/B CLKBUF1_27/Y NAND3X1_51/Y gnd vdd DFFPOSX1
XOAI21X1_79 INVX1_76/Y INVX1_79/Y AOI22X1_27/C gnd OAI21X1_80/C vdd OAI21X1
XNAND2X1_94 INVX1_76/A INVX1_79/Y gnd AOI22X1_26/D vdd NAND2X1
XAOI22X1_165 AOI22X1_165/A AND2X2_128/Y OAI21X1_499/C NOR2X1_220/Y gnd OAI21X1_502/C
+ vdd AOI22X1
XINVX1_345 INVX1_345/A gnd INVX1_345/Y vdd INVX1
XOAI21X1_524 INVX1_591/Y NAND2X1_502/Y OAI21X1_524/C gnd OAI21X1_524/Y vdd OAI21X1
XDFFPOSX1_163 INVX1_39/A CLKBUF1_38/Y OAI21X1_248/Y gnd vdd DFFPOSX1
XFILL_1_0_1 gnd vdd FILL
XFILL_19_1_2 gnd vdd FILL
XAOI22X1_72 NOR2X1_90/A INVX1_237/Y INVX1_239/Y AOI22X1_72/D gnd AOI22X1_72/Y vdd
+ AOI22X1
XDFFPOSX1_127 INVX1_207/A CLKBUF1_16/Y OAI21X1_193/Y gnd vdd DFFPOSX1
XNAND2X1_58 NAND2X1_58/A AOI22X1_13/Y gnd NAND2X1_58/Y vdd NAND2X1
XOAI21X1_43 NOR2X1_22/Y AOI21X1_4/Y BUFX2_143/A gnd NAND2X1_59/A vdd OAI21X1
XDFFPOSX1_61 INVX1_84/A CLKBUF1_3/Y NAND3X1_33/Y gnd vdd DFFPOSX1
XAOI22X1_129 NAND2X1_384/Y AND2X2_101/Y AOI22X1_129/C NOR2X1_166/Y gnd OAI21X1_394/C
+ vdd AOI22X1
XOAI21X1_488 INVX1_549/Y NAND2X1_469/Y OAI21X1_488/C gnd OAI21X1_488/Y vdd OAI21X1
XINVX1_309 BUFX2_70/Y gnd INVX1_309/Y vdd INVX1
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd BUFX2_88/A vdd NOR2X1
XFILL_8_2 gnd vdd FILL
XAOI22X1_36 AND2X2_4/B INVX1_111/Y NOR2X1_51/B AOI22X1_36/D gnd AOI22X1_36/Y vdd AOI22X1
XNAND2X1_22 NOR2X1_8/Y NOR2X1_11/Y gnd NOR2X1_12/A vdd NAND2X1
XDFFPOSX1_25 INVX1_36/A CLKBUF1_45/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XAOI21X1_1 AOI21X1_1/A INVX1_19/Y AOI21X1_1/C gnd AOI21X1_1/Y vdd AOI21X1
XINVX1_273 AND2X2_9/B gnd INVX1_273/Y vdd INVX1
XOAI21X1_452 INVX1_507/Y NAND2X1_436/Y OAI21X1_451/Y gnd OAI21X1_452/Y vdd OAI21X1
XNAND3X1_99 NAND3X1_99/A NAND3X1_98/Y NAND3X1_99/C gnd NAND3X1_99/Y vdd NAND3X1
XFILL_20_2_0 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XOAI21X1_416 INVX1_465/Y OAI21X1_416/B OAI21X1_416/C gnd OAI21X1_416/Y vdd OAI21X1
XNAND3X1_63 NOR2X1_74/Y NAND3X1_62/Y NAND3X1_63/C gnd NAND3X1_63/Y vdd NAND3X1
XNAND2X1_530 INVX1_623/A INVX1_624/A gnd NAND2X1_530/Y vdd NAND2X1
XFILL_26_1_2 gnd vdd FILL
XFILL_6_2_2 gnd vdd FILL
XFILL_8_0_1 gnd vdd FILL
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_201 BUFX2_31/Y gnd NOR2X1_78/B vdd INVX1
XOAI21X1_380 INVX1_423/Y OAI21X1_380/B OAI21X1_380/C gnd OAI21X1_380/Y vdd OAI21X1
XAND2X2_132 INVX1_606/A INVX1_599/A gnd AND2X2_132/Y vdd AND2X2
XNAND3X1_27 NOR2X1_35/Y NAND3X1_26/Y OAI21X1_66/Y gnd NAND3X1_27/Y vdd NAND3X1
XNAND2X1_494 INVX1_580/A INVX1_583/A gnd OAI21X1_518/B vdd NAND2X1
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XOAI21X1_344 INVX1_381/Y OAI21X1_344/B OAI21X1_343/Y gnd OAI21X1_344/Y vdd OAI21X1
XINVX1_47 INVX1_89/A gnd INVX1_47/Y vdd INVX1
XNAND2X1_458 BUFX2_62/Y INVX1_534/Y gnd NAND2X1_458/Y vdd NAND2X1
XAND2X2_69 INVX1_279/A INVX1_283/A gnd AND2X2_69/Y vdd AND2X2
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XFILL_7_3_0 gnd vdd FILL
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XFILL_27_2_0 gnd vdd FILL
XOAI21X1_308 INVX1_339/Y OAI21X1_308/B OAI21X1_308/C gnd OAI21X1_308/Y vdd OAI21X1
XNAND2X1_422 INVX1_485/A NAND2X1_421/Y gnd NAND2X1_422/Y vdd NAND2X1
XAND2X2_33 AND2X2_1/Y INVX1_66/A gnd AND2X2_33/Y vdd AND2X2
XOAI21X1_272 INVX1_294/Y OAI21X1_272/B NAND3X1_93/A gnd AOI21X1_43/C vdd OAI21X1
XNAND2X1_386 AND2X2_7/Y INVX1_440/Y gnd NAND2X1_386/Y vdd NAND2X1
XNOR2X1_72 gnd NOR2X1_72/B gnd NOR2X1_72/Y vdd NOR2X1
XOAI21X1_236 INVX1_256/Y AOI22X1_76/Y AOI22X1_77/Y gnd OAI21X1_236/Y vdd OAI21X1
XNAND2X1_350 INVX1_392/A BUFX2_36/Y gnd NAND2X1_350/Y vdd NAND2X1
XINVX1_598 AND2X2_99/B gnd INVX1_598/Y vdd INVX1
XNOR2X1_36 AND2X2_1/B INVX1_64/Y gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_182 BUFX2_9/Y INVX1_610/Y INVX1_611/Y gnd NAND3X1_183/B vdd NAND3X1
XNAND3X1_1 OR2X2_1/B INVX1_4/A NOR2X1_10/A gnd INVX1_2/A vdd NAND3X1
XOAI21X1_200 BUFX2_55/Y INVX1_218/Y INVX1_217/Y gnd OAI21X1_201/C vdd OAI21X1
XNOR2X1_233 gnd INVX1_586/Y gnd NOR2X1_233/Y vdd NOR2X1
XNAND2X1_314 BUFX2_84/Y INVX1_352/A gnd OAI21X1_320/B vdd NAND2X1
XNAND3X1_146 BUFX2_134/Y INVX1_484/Y INVX1_485/Y gnd NAND3X1_147/B vdd NAND3X1
XINVX1_562 INVX1_562/A gnd INVX1_562/Y vdd INVX1
XCLKBUF1_24 BUFX2_7/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOAI21X1_164 INVX1_167/A INVX1_174/Y OAI21X1_164/C gnd NAND3X1_59/C vdd OAI21X1
XNOR2X1_197 gnd INVX1_502/Y gnd NOR2X1_197/Y vdd NOR2X1
XNAND2X1_278 AND2X2_71/B NAND2X1_277/Y gnd AOI22X1_91/A vdd NAND2X1
XDFFPOSX1_344 INVX1_583/A CLKBUF1_47/Y AOI21X1_84/Y gnd vdd DFFPOSX1
XBUFX2_111 NOR3X1_4/Y gnd INVX1_421/A vdd BUFX2
XINVX1_526 INVX1_69/A gnd INVX1_526/Y vdd INVX1
XNAND3X1_110 BUFX2_122/Y INVX1_358/Y INVX1_359/Y gnd NAND3X1_110/Y vdd NAND3X1
XXNOR2X1_71 INVX1_69/A BUFX2_66/Y gnd AOI21X1_76/B vdd XNOR2X1
XOAI21X1_128 INVX1_132/Y INVX1_135/Y AOI22X1_43/C gnd OAI21X1_128/Y vdd OAI21X1
XNOR2X1_161 gnd INVX1_418/Y gnd NOR2X1_161/Y vdd NOR2X1
XNAND2X1_242 BUFX2_51/Y INVX1_261/Y gnd AOI22X1_78/D vdd NAND2X1
XDFFPOSX1_308 INVX1_520/A CLKBUF1_25/Y AOI21X1_75/Y gnd vdd DFFPOSX1
XINVX1_490 INVX1_490/A gnd INVX1_490/Y vdd INVX1
XXNOR2X1_35 BUFX2_58/Y AND2X2_9/Y gnd XNOR2X1_35/Y vdd XNOR2X1
XNOR2X1_125 gnd INVX1_334/Y gnd NOR2X1_125/Y vdd NOR2X1
XNAND2X1_206 BUFX2_55/Y INVX1_219/A gnd NAND2X1_206/Y vdd NAND2X1
XINVX1_454 BUFX2_114/Y gnd INVX1_454/Y vdd INVX1
XDFFPOSX1_272 AND2X2_9/A CLKBUF1_13/Y AOI21X1_66/Y gnd vdd DFFPOSX1
XNAND2X1_170 INVX1_168/A BUFX2_85/Y gnd NAND2X1_171/B vdd NAND2X1
XDFFPOSX1_236 INVX1_394/A CLKBUF1_44/Y AOI21X1_57/Y gnd vdd DFFPOSX1
XAOI21X1_68 INVX1_471/Y XNOR2X1_63/Y AOI21X1_68/C gnd AOI21X1_68/Y vdd AOI21X1
XINVX1_418 BUFX2_28/Y gnd INVX1_418/Y vdd INVX1
XBUFX2_71 BUFX2_67/A gnd INVX1_99/A vdd BUFX2
XNAND2X1_134 BUFX2_82/Y INVX1_125/Y gnd NAND2X1_134/Y vdd NAND2X1
XINVX1_382 AND2X2_88/B gnd INVX1_382/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XAOI21X1_32 INVX1_219/Y AOI21X1_32/B AOI21X1_32/C gnd AOI21X1_32/Y vdd AOI21X1
XDFFPOSX1_200 INVX1_331/A CLKBUF1_44/Y AOI21X1_48/Y gnd vdd DFFPOSX1
XBUFX2_35 RST_N gnd BUFX2_35/Y vdd BUFX2
XDFFPOSX1_98 AOI22X1_49/C CLKBUF1_15/Y OAI21X1_148/Y gnd vdd DFFPOSX1
XOAI21X1_80 INVX1_80/Y OAI21X1_80/B OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XNAND2X1_95 INVX1_77/A BUFX2_42/Y gnd NAND2X1_96/B vdd NAND2X1
XAOI22X1_166 INVX1_567/A INVX1_566/Y INVX1_568/Y NAND2X1_486/Y gnd OAI21X1_508/B vdd
+ AOI22X1
XINVX1_346 INVX1_88/A gnd INVX1_346/Y vdd INVX1
XOAI21X1_525 INVX1_588/Y OAI21X1_525/B NOR2X1_233/Y gnd AOI21X1_85/C vdd OAI21X1
XDFFPOSX1_164 INVX1_268/A CLKBUF1_46/Y AOI21X1_39/Y gnd vdd DFFPOSX1
XFILL_1_0_2 gnd vdd FILL
XAOI22X1_73 AOI22X1_73/A AND2X2_62/Y AOI22X1_73/C NOR2X1_90/Y gnd AOI22X1_73/Y vdd
+ AOI22X1
XNAND2X1_59 NAND2X1_59/A AOI22X1_14/Y gnd NAND2X1_59/Y vdd NAND2X1
XDFFPOSX1_128 INVX1_205/A CLKBUF1_16/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_62 AOI22X1_31/C CLKBUF1_3/Y OAI21X1_92/Y gnd vdd DFFPOSX1
XOAI21X1_44 NOR2X1_24/Y AND2X2_25/Y INVX1_38/A gnd AND2X2_26/B vdd OAI21X1
XAOI22X1_130 INVX1_441/A INVX1_440/Y INVX1_442/Y AOI22X1_130/D gnd OAI21X1_400/B vdd
+ AOI22X1
XOAI21X1_489 INVX1_546/Y NAND2X1_470/Y NOR2X1_215/Y gnd AOI21X1_79/C vdd OAI21X1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XAOI22X1_37 AOI22X1_37/A AND2X2_41/Y AOI22X1_37/C NOR2X1_51/Y gnd AOI22X1_37/Y vdd
+ AOI22X1
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd BUFX2_96/A vdd NOR2X1
XFILL_8_3 gnd vdd FILL
XDFFPOSX1_26 INVX1_37/A CLKBUF1_20/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XNAND2X1_23 INVX1_5/A BUFX2_70/Y gnd NAND2X1_23/Y vdd NAND2X1
XINVX1_274 BUFX2_58/Y gnd INVX1_274/Y vdd INVX1
XAOI21X1_2 INVX1_19/Y EN_request_put INVX1_3/Y gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_453 INVX1_504/Y NAND2X1_437/Y NOR2X1_197/Y gnd AOI21X1_73/C vdd OAI21X1
XFILL_22_0_0 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XFILL_20_2_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XINVX1_238 NOR2X1_90/A gnd INVX1_238/Y vdd INVX1
XOAI21X1_417 INVX1_462/Y OAI21X1_417/B NOR2X1_179/Y gnd AOI21X1_67/C vdd OAI21X1
XNAND3X1_64 AND2X2_8/Y NOR2X1_77/B INVX1_198/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND2X1_531 AND2X2_21/A NAND2X1_530/Y gnd NAND2X1_531/Y vdd NAND2X1
XFILL_8_0_2 gnd vdd FILL
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_202 INVX1_484/A gnd INVX1_202/Y vdd INVX1
XOAI21X1_381 INVX1_420/Y OAI21X1_381/B NOR2X1_161/Y gnd AOI21X1_61/C vdd OAI21X1
XNAND3X1_28 INVX1_69/A INVX1_71/Y INVX1_72/Y gnd NAND3X1_29/B vdd NAND3X1
XAND2X2_133 INVX1_606/A INVX1_592/A gnd NOR2X1_230/B vdd AND2X2
XNAND2X1_495 INVX1_582/A INVX1_580/Y gnd NAND2X1_495/Y vdd NAND2X1
XINVX1_166 BUFX2_34/Y gnd INVX1_166/Y vdd INVX1
XOAI21X1_345 INVX1_378/Y OAI21X1_345/B NOR2X1_143/Y gnd AOI21X1_55/C vdd OAI21X1
XINVX1_48 BUFX2_56/Y gnd INVX1_48/Y vdd INVX1
XFILL_12_1 gnd vdd FILL
XNAND2X1_459 INVX1_532/A INVX1_244/A gnd NAND2X1_460/B vdd NAND2X1
XAND2X2_70 INVX1_575/A INVX1_578/A gnd AND2X2_70/Y vdd AND2X2
XFILL_27_2_1 gnd vdd FILL
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XFILL_7_3_1 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XINVX1_130 AND2X2_99/B gnd INVX1_130/Y vdd INVX1
XOAI21X1_309 INVX1_336/Y NAND2X1_305/Y NOR2X1_125/Y gnd AOI21X1_49/C vdd OAI21X1
XNAND2X1_423 INVX1_463/A AND2X2_11/A gnd NAND2X1_423/Y vdd NAND2X1
XAND2X2_34 INVX1_69/A INVX1_73/A gnd AND2X2_34/Y vdd AND2X2
XNAND2X1_387 INVX1_440/A INVX1_443/Y gnd AOI22X1_130/D vdd NAND2X1
XOAI21X1_273 INVX1_298/Y AOI22X1_88/Y AOI22X1_89/Y gnd OAI21X1_273/Y vdd OAI21X1
XNOR2X1_73 NOR2X1_73/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XOAI21X1_237 BUFX2_51/Y INVX1_260/Y INVX1_259/Y gnd OAI21X1_237/Y vdd OAI21X1
XNAND2X1_351 INVX1_394/A NAND2X1_350/Y gnd NAND2X1_351/Y vdd NAND2X1
XNAND3X1_183 NOR2X1_239/Y NAND3X1_183/B NAND3X1_183/C gnd NAND3X1_183/Y vdd NAND3X1
XINVX1_599 INVX1_599/A gnd INVX1_599/Y vdd INVX1
XNOR2X1_37 gnd INVX1_68/Y gnd NOR2X1_37/Y vdd NOR2X1
XNAND3X1_2 INVX1_1/Y INVX1_2/Y NOR2X1_8/Y gnd INVX1_3/A vdd NAND3X1
XOAI21X1_201 INVX1_209/A INVX1_216/Y OAI21X1_201/C gnd NAND3X1_71/C vdd OAI21X1
XNOR2X1_234 INVX1_588/A INVX1_589/Y gnd NOR2X1_234/Y vdd NOR2X1
XNAND2X1_315 BUFX2_118/Y INVX1_349/Y gnd NAND2X1_315/Y vdd NAND2X1
XNAND3X1_147 NOR2X1_185/Y NAND3X1_147/B OAI21X1_432/Y gnd NAND3X1_147/Y vdd NAND3X1
XINVX1_563 INVX1_479/A gnd INVX1_563/Y vdd INVX1
XCLKBUF1_25 BUFX2_2/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XOR2X2_5 OR2X2_5/A OR2X2_4/B gnd OR2X2_5/Y vdd OR2X2
XOAI21X1_165 INVX1_174/Y INVX1_177/Y AOI22X1_55/C gnd OAI21X1_166/C vdd OAI21X1
XNOR2X1_198 NAND2X1_2/B INVX1_505/Y gnd NOR2X1_198/Y vdd NOR2X1
XNAND2X1_279 BUFX2_21/Y INVX1_310/A gnd NAND2X1_279/Y vdd NAND2X1
XDFFPOSX1_345 INVX1_581/A CLKBUF1_47/Y NAND3X1_175/Y gnd vdd DFFPOSX1
XBUFX2_112 NOR3X1_4/Y gnd BUFX2_112/Y vdd BUFX2
XINVX1_527 AND2X2_13/A gnd INVX1_527/Y vdd INVX1
XNAND3X1_111 NOR2X1_131/Y NAND3X1_110/Y OAI21X1_324/Y gnd NAND3X1_111/Y vdd NAND3X1
XNOR2X1_162 INVX1_420/A INVX1_421/Y gnd NOR2X1_162/Y vdd NOR2X1
XOAI21X1_129 INVX1_136/Y NAND2X1_138/Y OAI21X1_128/Y gnd OAI21X1_129/Y vdd OAI21X1
XXNOR2X1_72 INVX1_244/A BUFX2_62/Y gnd XNOR2X1_72/Y vdd XNOR2X1
XNAND2X1_243 NOR2X1_97/A INVX1_251/A gnd NAND2X1_243/Y vdd NAND2X1
XINVX1_491 INVX1_237/A gnd INVX1_491/Y vdd INVX1
XDFFPOSX1_309 INVX1_518/A CLKBUF1_29/Y NAND3X1_157/Y gnd vdd DFFPOSX1
XXNOR2X1_36 BUFX2_57/Y INVX1_279/A gnd AOI21X1_41/B vdd XNOR2X1
XNAND2X1_207 INVX1_209/A INVX1_216/Y gnd OAI21X1_204/B vdd NAND2X1
XNOR2X1_126 INVX1_336/A INVX1_337/Y gnd NOR2X1_126/Y vdd NOR2X1
XDFFPOSX1_273 INVX1_455/A CLKBUF1_13/Y NAND3X1_139/Y gnd vdd DFFPOSX1
XINVX1_455 INVX1_455/A gnd INVX1_455/Y vdd INVX1
XNAND2X1_171 INVX1_170/A NAND2X1_171/B gnd AOI22X1_53/A vdd NAND2X1
XAOI21X1_69 INVX1_478/Y XNOR2X1_64/Y AOI21X1_69/C gnd AOI21X1_69/Y vdd AOI21X1
XDFFPOSX1_237 INVX1_392/A CLKBUF1_7/Y NAND3X1_121/Y gnd vdd DFFPOSX1
XINVX1_419 BUFX2_80/Y gnd INVX1_419/Y vdd INVX1
XBUFX2_72 BUFX2_67/A gnd BUFX2_72/Y vdd BUFX2
XFILL_15_0_1 gnd vdd FILL
XNAND2X1_135 INVX1_125/A INVX1_128/Y gnd AOI22X1_40/D vdd NAND2X1
XAOI21X1_33 INVX1_226/Y XNOR2X1_28/Y AOI21X1_33/C gnd AOI21X1_33/Y vdd AOI21X1
XFILL_13_2_2 gnd vdd FILL
XINVX1_383 INVX1_96/A gnd INVX1_383/Y vdd INVX1
XDFFPOSX1_201 AND2X2_21/B CLKBUF1_7/Y NAND3X1_103/Y gnd vdd DFFPOSX1
XBUFX2_36 BUFX2_39/A gnd BUFX2_36/Y vdd BUFX2
XDFFPOSX1_99 INVX1_158/A CLKBUF1_15/Y DFFPOSX1_99/D gnd vdd DFFPOSX1
XNAND2X1_96 INVX1_79/A NAND2X1_96/B gnd AOI22X1_27/A vdd NAND2X1
XOAI21X1_81 INVX1_77/Y OAI21X1_81/B NOR2X1_39/Y gnd OAI21X1_81/Y vdd OAI21X1
XDFFPOSX1_165 NOR2X1_99/A CLKBUF1_46/Y NAND3X1_85/Y gnd vdd DFFPOSX1
XAOI22X1_167 AOI22X1_167/A AND2X2_129/Y AOI22X1_167/C NOR2X1_222/Y gnd OAI21X1_508/C
+ vdd AOI22X1
XINVX1_347 AND2X2_80/A gnd INVX1_347/Y vdd INVX1
XOAI21X1_526 INVX1_592/Y OAI21X1_526/B OAI21X1_526/C gnd OAI21X1_526/Y vdd OAI21X1
XAOI22X1_74 INVX1_245/A INVX1_244/Y NOR2X1_92/B AOI22X1_74/D gnd AOI22X1_74/Y vdd
+ AOI22X1
XNAND2X1_60 OR2X2_5/A OR2X2_3/B gnd AOI21X1_5/B vdd NAND2X1
XOAI21X1_45 NOR2X1_25/Y AND2X2_27/Y INVX1_39/Y gnd OAI21X1_45/Y vdd OAI21X1
XDFFPOSX1_129 AND2X2_10/B CLKBUF1_16/Y NAND3X1_67/Y gnd vdd DFFPOSX1
XAOI22X1_131 NAND2X1_389/Y AND2X2_102/Y OAI21X1_397/C NOR2X1_168/Y gnd OAI21X1_400/C
+ vdd AOI22X1
XDFFPOSX1_63 INVX1_87/A CLKBUF1_7/Y OAI21X1_94/Y gnd vdd DFFPOSX1
XINVX1_311 AND2X2_74/B gnd INVX1_311/Y vdd INVX1
XFILL_14_3_0 gnd vdd FILL
XOAI21X1_490 INVX1_550/Y OAI21X1_490/B AOI22X1_161/Y gnd OAI21X1_490/Y vdd OAI21X1
XAOI22X1_38 NOR2X1_53/A INVX1_118/Y NOR2X1_53/B AOI22X1_38/D gnd AOI22X1_38/Y vdd
+ AOI22X1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd BUFX2_98/A vdd NOR2X1
XDFFPOSX1_27 BUFX2_137/A CLKBUF1_20/Y NAND2X1_53/Y gnd vdd DFFPOSX1
XNAND2X1_24 INVX1_3/A NAND2X1_23/Y gnd BUFX2_54/A vdd NAND2X1
XAOI21X1_3 AND2X2_24/Y INVX1_31/Y AOI21X1_3/C gnd AOI21X1_3/Y vdd AOI21X1
XINVX1_275 INVX1_275/A gnd INVX1_275/Y vdd INVX1
XOAI21X1_454 INVX1_508/Y AOI22X1_148/Y AOI22X1_149/Y gnd OAI21X1_454/Y vdd OAI21X1
XFILL_22_0_1 gnd vdd FILL
XFILL_0_3_2 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XFILL_20_2_2 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XINVX1_239 BUFX2_17/Y gnd INVX1_239/Y vdd INVX1
XOAI21X1_418 INVX1_466/Y AOI22X1_136/Y AOI22X1_137/Y gnd OAI21X1_418/Y vdd OAI21X1
XNAND3X1_65 NOR2X1_76/Y NAND3X1_64/Y NAND3X1_65/C gnd NAND3X1_65/Y vdd NAND3X1
XINVX1_203 AND2X2_10/B gnd INVX1_203/Y vdd INVX1
XOAI21X1_382 INVX1_424/Y OAI21X1_382/B OAI21X1_382/C gnd OAI21X1_382/Y vdd OAI21X1
XINVX1_85 BUFX2_76/Y gnd INVX1_85/Y vdd INVX1
XNAND3X1_29 NOR2X1_37/Y NAND3X1_29/B OAI21X1_72/Y gnd NAND3X1_29/Y vdd NAND3X1
XAND2X2_134 INVX1_599/A INVX1_592/A gnd AND2X2_134/Y vdd AND2X2
XNAND2X1_496 INVX1_580/A INVX1_583/Y gnd AOI22X1_170/D vdd NAND2X1
XINVX1_49 INVX1_4/A gnd INVX1_49/Y vdd INVX1
XFILL_21_3_0 gnd vdd FILL
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XOAI21X1_346 INVX1_382/Y OAI21X1_346/B OAI21X1_346/C gnd OAI21X1_346/Y vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XNAND2X1_460 AND2X2_14/A NAND2X1_460/B gnd NAND2X1_460/Y vdd NAND2X1
XAND2X2_71 INVX1_294/A AND2X2_71/B gnd INVX1_293/A vdd AND2X2
XFILL_9_1_1 gnd vdd FILL
XFILL_27_2_2 gnd vdd FILL
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XFILL_7_3_2 gnd vdd FILL
XINVX1_131 INVX1_89/A gnd NOR2X1_57/B vdd INVX1
XOAI21X1_310 INVX1_340/Y AOI22X1_100/Y OAI21X1_310/C gnd OAI21X1_310/Y vdd OAI21X1
XNAND2X1_424 INVX1_237/A INVX1_489/Y gnd OAI21X1_441/B vdd NAND2X1
XAND2X2_35 INVX1_76/A INVX1_80/A gnd AND2X2_35/Y vdd AND2X2
XOAI21X1_274 BUFX2_52/Y INVX1_302/Y INVX1_301/Y gnd OAI21X1_274/Y vdd OAI21X1
XNAND2X1_388 INVX1_441/A AND2X2_7/Y gnd NAND2X1_389/B vdd NAND2X1
XNOR2X1_74 gnd NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XFILL_28_3_0 gnd vdd FILL
XOAI21X1_238 INVX1_251/A INVX1_258/Y OAI21X1_237/Y gnd NAND3X1_83/C vdd OAI21X1
XNAND2X1_352 BUFX2_38/Y AND2X2_4/A gnd OAI21X1_362/B vdd NAND2X1
XNAND3X1_184 BUFX2_8/Y INVX1_617/Y INVX1_618/Y gnd NAND3X1_185/B vdd NAND3X1
XINVX1_600 INVX1_96/A gnd INVX1_600/Y vdd INVX1
XNOR2X1_38 INVX1_70/A INVX1_71/Y gnd NOR2X1_38/Y vdd NOR2X1
XNAND3X1_3 INVX1_1/Y NAND3X1_3/B NOR2X1_9/Y gnd NOR2X1_12/B vdd NAND3X1
XNAND2X1_316 BUFX2_86/Y INVX1_352/Y gnd AOI22X1_104/D vdd NAND2X1
XOAI21X1_202 INVX1_216/Y INVX1_219/Y AOI22X1_67/C gnd OAI21X1_202/Y vdd OAI21X1
XNOR2X1_235 gnd INVX1_593/Y gnd NOR2X1_235/Y vdd NOR2X1
XNAND3X1_148 BUFX2_129/Y INVX1_491/Y INVX1_492/Y gnd NAND3X1_148/Y vdd NAND3X1
XINVX1_564 INVX1_564/A gnd INVX1_564/Y vdd INVX1
XCLKBUF1_26 BUFX2_4/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XOAI21X1_166 INVX1_178/Y OAI21X1_166/B OAI21X1_166/C gnd OAI21X1_166/Y vdd OAI21X1
XNOR2X1_199 gnd INVX1_509/Y gnd NOR2X1_199/Y vdd NOR2X1
XNAND2X1_280 INVX1_99/A INVX1_307/Y gnd NAND2X1_280/Y vdd NAND2X1
XNAND3X1_112 INVX1_363/A INVX1_365/Y INVX1_366/Y gnd NAND3X1_112/Y vdd NAND3X1
XDFFPOSX1_346 AOI22X1_173/C CLKBUF1_2/Y OAI21X1_524/Y gnd vdd DFFPOSX1
XBUFX2_113 NOR3X1_4/Y gnd BUFX2_113/Y vdd BUFX2
XINVX1_528 INVX1_528/A gnd INVX1_528/Y vdd INVX1
XNOR2X1_163 gnd INVX1_425/Y gnd NOR2X1_163/Y vdd NOR2X1
XXNOR2X1_73 INVX1_279/A BUFX2_64/Y gnd AOI21X1_78/B vdd XNOR2X1
XOAI21X1_130 INVX1_133/Y NAND2X1_139/Y NOR2X1_57/Y gnd AOI21X1_20/C vdd OAI21X1
XNAND2X1_244 AND2X2_64/B NAND2X1_243/Y gnd AOI22X1_79/A vdd NAND2X1
XINVX1_492 AND2X2_11/A gnd INVX1_492/Y vdd INVX1
XDFFPOSX1_310 AOI22X1_155/C CLKBUF1_21/Y OAI21X1_470/Y gnd vdd DFFPOSX1
XXNOR2X1_37 BUFX2_57/Y INVX1_575/A gnd AOI21X1_42/B vdd XNOR2X1
XNAND2X1_208 BUFX2_55/Y INVX1_219/Y gnd AOI22X1_66/D vdd NAND2X1
XNOR2X1_127 gnd INVX1_341/Y gnd NOR2X1_127/Y vdd NOR2X1
XDFFPOSX1_274 AOI22X1_137/C CLKBUF1_36/Y OAI21X1_416/Y gnd vdd DFFPOSX1
XINVX1_456 AND2X2_9/Y gnd INVX1_456/Y vdd INVX1
XNAND2X1_172 BUFX2_54/Y AND2X2_50/B gnd OAI21X1_166/B vdd NAND2X1
XAOI21X1_70 INVX1_485/Y AOI21X1_70/B AOI21X1_70/C gnd AOI21X1_70/Y vdd AOI21X1
XDFFPOSX1_238 OAI21X1_361/C CLKBUF1_39/Y OAI21X1_362/Y gnd vdd DFFPOSX1
XINVX1_420 INVX1_420/A gnd INVX1_420/Y vdd INVX1
XBUFX2_73 BUFX2_73/A gnd BUFX2_73/Y vdd BUFX2
XFILL_15_0_2 gnd vdd FILL
XNAND2X1_136 NOR2X1_56/A BUFX2_82/Y gnd NAND2X1_137/B vdd NAND2X1
XAOI21X1_34 INVX1_233/Y XNOR2X1_29/Y AOI21X1_34/C gnd AOI21X1_34/Y vdd AOI21X1
XINVX1_384 BUFX2_81/Y gnd INVX1_384/Y vdd INVX1
XDFFPOSX1_202 OAI21X1_307/C CLKBUF1_14/Y OAI21X1_308/Y gnd vdd DFFPOSX1
XBUFX2_37 BUFX2_39/A gnd BUFX2_37/Y vdd BUFX2
XNAND2X1_97 INVX1_114/A INVX1_107/A gnd NOR2X1_41/A vdd NAND2X1
XNAND2X1_100 BUFX2_76/Y INVX1_83/Y gnd OAI21X1_87/B vdd NAND2X1
XDFFPOSX1_166 AOI22X1_83/C CLKBUF1_20/Y OAI21X1_253/Y gnd vdd DFFPOSX1
XOAI21X1_82 INVX1_81/Y OAI21X1_82/B AOI22X1_27/Y gnd OAI21X1_82/Y vdd OAI21X1
XAOI22X1_168 INVX1_574/A INVX1_573/Y INVX1_575/Y NAND2X1_491/Y gnd AOI22X1_168/Y vdd
+ AOI22X1
XINVX1_348 BUFX2_28/Y gnd INVX1_348/Y vdd INVX1
XOAI21X1_527 BUFX2_78/Y INVX1_596/Y INVX1_595/Y gnd OAI21X1_528/C vdd OAI21X1
XAOI22X1_75 AOI22X1_75/A AND2X2_63/Y AOI22X1_75/C NOR2X1_92/Y gnd AOI22X1_75/Y vdd
+ AOI22X1
XDFFPOSX1_64 INVX1_93/A CLKBUF1_3/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XOAI21X1_46 INVX1_41/A INVX1_43/Y INVX1_42/Y gnd OAI21X1_47/C vdd OAI21X1
XFILL_25_1 gnd vdd FILL
XNAND2X1_61 OR2X2_4/A OR2X2_4/B gnd NAND2X1_61/Y vdd NAND2X1
XAOI22X1_132 INVX1_448/A INVX1_447/Y INVX1_449/Y AOI22X1_132/D gnd OAI21X1_406/B vdd
+ AOI22X1
XOAI21X1_491 BUFX2_97/Y INVX1_554/Y INVX1_553/Y gnd OAI21X1_491/Y vdd OAI21X1
XFILL_16_1_0 gnd vdd FILL
XDFFPOSX1_130 AOI22X1_65/C CLKBUF1_34/Y OAI21X1_197/Y gnd vdd DFFPOSX1
XINVX1_312 INVX1_38/A gnd INVX1_312/Y vdd INVX1
XFILL_14_3_1 gnd vdd FILL
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI22X1_39 AOI22X1_39/A AND2X2_42/Y AOI22X1_39/C NOR2X1_53/Y gnd AOI22X1_39/Y vdd
+ AOI22X1
XDFFPOSX1_28 BUFX2_138/A CLKBUF1_6/Y NAND2X1_54/Y gnd vdd DFFPOSX1
XOAI21X1_10 INVX1_18/Y NOR2X1_17/Y NAND2X1_29/Y gnd OAI21X1_10/Y vdd OAI21X1
XNAND2X1_25 NOR2X1_13/Y NOR2X1_14/Y gnd NOR3X1_1/B vdd NAND2X1
XAOI21X1_4 INVX1_31/Y INVX1_27/A EN_response_get gnd AOI21X1_4/Y vdd AOI21X1
XINVX1_276 INVX1_459/A gnd INVX1_276/Y vdd INVX1
XOAI21X1_455 BUFX2_89/Y INVX1_512/Y INVX1_511/Y gnd OAI21X1_455/Y vdd OAI21X1
XFILL_22_0_2 gnd vdd FILL
XFILL_2_1_2 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XNAND3X1_66 INVX1_484/A NOR2X1_79/B INVX1_205/Y gnd NAND3X1_66/Y vdd NAND3X1
XOAI21X1_419 BUFX2_90/Y INVX1_470/Y INVX1_469/Y gnd OAI21X1_419/Y vdd OAI21X1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XINVX1_204 INVX1_204/A gnd NOR2X1_79/B vdd INVX1
XOAI21X1_383 BUFX2_87/Y INVX1_428/Y INVX1_427/Y gnd OAI21X1_383/Y vdd OAI21X1
XAND2X2_135 BUFX2_26/Y INVX1_46/A gnd AND2X2_135/Y vdd AND2X2
XNAND3X1_30 INVX1_76/A INVX1_78/Y INVX1_79/Y gnd NAND3X1_30/Y vdd NAND3X1
XNAND2X1_497 INVX1_581/A INVX1_582/A gnd NAND2X1_498/B vdd NAND2X1
XFILL_23_1_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XINVX1_50 INVX1_41/A gnd INVX1_50/Y vdd INVX1
XFILL_21_3_1 gnd vdd FILL
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XOAI21X1_347 BUFX2_81/Y INVX1_386/Y INVX1_385/Y gnd OAI21X1_347/Y vdd OAI21X1
XFILL_12_3 gnd vdd FILL
XNAND2X1_461 BUFX2_64/Y AND2X2_15/A gnd OAI21X1_482/B vdd NAND2X1
XAND2X2_72 INVX1_293/A AND2X2_72/B gnd AND2X2_72/Y vdd AND2X2
XFILL_9_1_2 gnd vdd FILL
XOAI21X1_311 BUFX2_77/Y INVX1_344/Y INVX1_343/Y gnd OAI21X1_311/Y vdd OAI21X1
XINVX1_14 BUFX2_30/Y gnd INVX1_14/Y vdd INVX1
XINVX1_132 BUFX2_50/Y gnd INVX1_132/Y vdd INVX1
XNAND2X1_425 BUFX2_129/Y INVX1_492/Y gnd AOI22X1_144/D vdd NAND2X1
XAND2X2_36 INVX1_84/A INVX1_93/A gnd INVX1_83/A vdd AND2X2
XOAI21X1_275 INVX1_293/A INVX1_300/Y OAI21X1_274/Y gnd NAND3X1_95/C vdd OAI21X1
XNAND2X1_389 AND2X2_7/A NAND2X1_389/B gnd NAND2X1_389/Y vdd NAND2X1
XNOR2X1_75 AND2X2_3/B NOR2X1_75/B gnd NOR2X1_75/Y vdd NOR2X1
XFILL_28_3_1 gnd vdd FILL
XOAI21X1_239 INVX1_258/Y INVX1_261/Y AOI22X1_79/C gnd OAI21X1_239/Y vdd OAI21X1
XNAND2X1_353 AND2X2_4/Y INVX1_398/Y gnd OAI21X1_363/B vdd NAND2X1
XNAND3X1_185 NOR2X1_241/Y NAND3X1_185/B OAI21X1_546/Y gnd NAND3X1_185/Y vdd NAND3X1
XINVX1_601 INVX1_601/A gnd INVX1_601/Y vdd INVX1
XNAND3X1_4 INVX1_7/Y NAND3X1_3/B NOR2X1_8/Y gnd NOR3X1_1/C vdd NAND3X1
XOAI21X1_203 INVX1_220/Y NAND2X1_206/Y OAI21X1_202/Y gnd OAI21X1_203/Y vdd OAI21X1
XNOR2X1_39 gnd INVX1_75/Y gnd NOR2X1_39/Y vdd NOR2X1
XNAND2X1_317 NAND2X1_7/A BUFX2_118/Y gnd NAND2X1_317/Y vdd NAND2X1
XNOR2X1_236 NAND2X1_6/B INVX1_596/Y gnd NOR2X1_236/Y vdd NOR2X1
XCLKBUF1_27 BUFX2_1/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XNAND3X1_149 NOR2X1_187/Y NAND3X1_148/Y OAI21X1_438/Y gnd NAND3X1_149/Y vdd NAND3X1
XINVX1_565 BUFX2_28/Y gnd INVX1_565/Y vdd INVX1
XOAI21X1_167 INVX1_175/Y NAND2X1_173/Y NOR2X1_70/Y gnd AOI21X1_26/C vdd OAI21X1
XNOR2X1_200 INVX1_511/A INVX1_512/Y gnd NOR2X1_200/Y vdd NOR2X1
XNAND2X1_281 BUFX2_21/Y INVX1_310/Y gnd AOI22X1_92/D vdd NAND2X1
XNAND3X1_113 NOR2X1_133/Y NAND3X1_112/Y NAND3X1_113/C gnd NAND3X1_113/Y vdd NAND3X1
XBUFX2_114 NOR3X1_4/Y gnd BUFX2_114/Y vdd BUFX2
XINVX1_529 INVX1_73/A gnd INVX1_529/Y vdd INVX1
XDFFPOSX1_347 INVX1_592/A CLKBUF1_14/Y OAI21X1_526/Y gnd vdd DFFPOSX1
XXNOR2X1_74 INVX1_547/A BUFX2_74/Y gnd AOI21X1_79/B vdd XNOR2X1
XNOR2X1_164 INVX1_427/A INVX1_428/Y gnd NOR2X1_164/Y vdd NOR2X1
XOAI21X1_131 INVX1_137/Y AOI22X1_42/Y AOI22X1_43/Y gnd DFFPOSX1_87/D vdd OAI21X1
XNAND2X1_245 BUFX2_60/Y INVX1_268/A gnd NAND2X1_245/Y vdd NAND2X1
XDFFPOSX1_311 INVX1_73/A CLKBUF1_51/Y OAI21X1_472/Y gnd vdd DFFPOSX1
XINVX1_493 INVX1_493/A gnd INVX1_493/Y vdd INVX1
XXNOR2X1_38 BUFX2_100/Y INVX1_293/A gnd AOI21X1_43/B vdd XNOR2X1
XNOR2X1_128 INVX1_343/A INVX1_344/Y gnd NOR2X1_128/Y vdd NOR2X1
XNAND2X1_209 INVX1_217/A INVX1_209/A gnd NAND2X1_210/B vdd NAND2X1
XDFFPOSX1_275 INVX1_466/A CLKBUF1_42/Y OAI21X1_418/Y gnd vdd DFFPOSX1
XINVX1_457 AND2X2_9/A gnd INVX1_457/Y vdd INVX1
XNAND2X1_173 INVX1_167/A INVX1_174/Y gnd NAND2X1_173/Y vdd NAND2X1
XAOI21X1_71 INVX1_492/Y XNOR2X1_66/Y AOI21X1_71/C gnd AOI21X1_71/Y vdd AOI21X1
XINVX1_421 INVX1_421/A gnd INVX1_421/Y vdd INVX1
XDFFPOSX1_239 INVX1_115/A CLKBUF1_39/Y OAI21X1_364/Y gnd vdd DFFPOSX1
XBUFX2_74 BUFX2_73/A gnd BUFX2_74/Y vdd BUFX2
XNAND2X1_137 NAND2X1_5/B NAND2X1_137/B gnd AOI22X1_41/A vdd NAND2X1
XAOI21X1_35 INVX1_240/Y XNOR2X1_30/Y AOI21X1_35/C gnd AOI21X1_35/Y vdd AOI21X1
XDFFPOSX1_203 AND2X2_79/B CLKBUF1_14/Y OAI21X1_310/Y gnd vdd DFFPOSX1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XBUFX2_38 BUFX2_39/A gnd BUFX2_38/Y vdd BUFX2
XNAND2X1_98 INVX1_98/A INVX1_121/A gnd NOR2X1_41/B vdd NAND2X1
XOAI21X1_83 INVX1_83/A INVX1_85/Y INVX1_84/Y gnd OAI21X1_83/Y vdd OAI21X1
XNAND2X1_101 INVX1_83/A INVX1_86/Y gnd AOI22X1_28/D vdd NAND2X1
XINVX1_349 BUFX2_86/Y gnd INVX1_349/Y vdd INVX1
XDFFPOSX1_167 INVX1_277/A CLKBUF1_28/Y OAI21X1_255/Y gnd vdd DFFPOSX1
XAOI22X1_169 AOI22X1_169/A AND2X2_130/Y AOI22X1_169/C NOR2X1_224/Y gnd AOI22X1_169/Y
+ vdd AOI22X1
XFILL_3_1 gnd vdd FILL
XOAI21X1_528 BUFX2_13/Y INVX1_594/Y OAI21X1_528/C gnd NAND3X1_179/C vdd OAI21X1
XAOI22X1_76 NOR2X1_95/A INVX1_251/Y INVX1_253/Y AOI22X1_76/D gnd AOI22X1_76/Y vdd
+ AOI22X1
XDFFPOSX1_65 INVX1_91/A CLKBUF1_12/Y NAND3X1_35/Y gnd vdd DFFPOSX1
XOAI21X1_47 BUFX2_24/Y INVX1_41/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XFILL_25_2 gnd vdd FILL
XNAND2X1_62 OR2X2_5/A OR2X2_4/B gnd NAND3X1_19/B vdd NAND2X1
XAOI22X1_133 AOI22X1_133/A AND2X2_103/Y AOI22X1_133/C NOR2X1_170/Y gnd OAI21X1_406/C
+ vdd AOI22X1
XOAI21X1_492 INVX1_554/A INVX1_552/Y OAI21X1_491/Y gnd OAI21X1_492/Y vdd OAI21X1
XFILL_16_1_1 gnd vdd FILL
XDFFPOSX1_131 INVX1_395/A CLKBUF1_5/Y OAI21X1_199/Y gnd vdd DFFPOSX1
XINVX1_313 BUFX2_30/Y gnd INVX1_313/Y vdd INVX1
XFILL_14_3_2 gnd vdd FILL
XNOR2X1_9 INVX1_7/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI22X1_40 NOR2X1_56/A INVX1_125/Y NOR2X1_56/B AOI22X1_40/D gnd AOI22X1_40/Y vdd
+ AOI22X1
XNAND2X1_26 NOR2X1_10/A INVX1_3/A gnd NAND2X1_26/Y vdd NAND2X1
XDFFPOSX1_29 BUFX2_139/A CLKBUF1_6/Y NAND2X1_55/Y gnd vdd DFFPOSX1
XOAI21X1_11 INVX1_20/Y NOR2X1_17/Y OAI21X1_11/C gnd DFFPOSX1_5/D vdd OAI21X1
XINVX1_277 INVX1_277/A gnd INVX1_277/Y vdd INVX1
XOAI21X1_456 BUFX2_63/Y INVX1_510/Y OAI21X1_455/Y gnd OAI21X1_456/Y vdd OAI21X1
XAOI21X1_5 OR2X2_3/Y AOI21X1_5/B INVX1_38/Y gnd AOI21X1_6/C vdd AOI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XOAI21X1_420 BUFX2_132/Y INVX1_468/Y OAI21X1_419/Y gnd OAI21X1_420/Y vdd OAI21X1
XNAND3X1_67 NOR2X1_78/Y NAND3X1_66/Y NAND3X1_67/C gnd NAND3X1_67/Y vdd NAND3X1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XOAI21X1_384 BUFX2_116/Y INVX1_426/Y OAI21X1_383/Y gnd OAI21X1_384/Y vdd OAI21X1
XAND2X2_136 BUFX2_81/Y AND2X2_99/B gnd AND2X2_136/Y vdd AND2X2
XNAND3X1_31 NOR2X1_39/Y NAND3X1_30/Y OAI21X1_78/Y gnd NAND3X1_31/Y vdd NAND3X1
XNAND2X1_498 INVX1_583/A NAND2X1_498/B gnd AOI22X1_171/A vdd NAND2X1
XFILL_5_0_0 gnd vdd FILL
XFILL_23_1_1 gnd vdd FILL
XFILL_21_3_2 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_169 BUFX2_85/Y gnd INVX1_169/Y vdd INVX1
XAND2X2_100 BUFX2_84/Y INVX1_430/A gnd AND2X2_100/Y vdd AND2X2
XOAI21X1_348 BUFX2_37/Y INVX1_384/Y OAI21X1_347/Y gnd NAND3X1_119/C vdd OAI21X1
XNAND2X1_462 INVX1_279/A INVX1_538/Y gnd NAND2X1_462/Y vdd NAND2X1
XAND2X2_73 BUFX2_51/Y AND2X2_73/B gnd AND2X2_73/Y vdd AND2X2
XINVX1_15 EN_request_put gnd INVX1_15/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XOAI21X1_312 AND2X2_85/A INVX1_342/Y OAI21X1_311/Y gnd NAND3X1_107/C vdd OAI21X1
XNAND2X1_426 INVX1_490/A INVX1_237/A gnd NAND2X1_427/B vdd NAND2X1
XAND2X2_37 INVX1_83/A INVX1_87/A gnd AND2X2_37/Y vdd AND2X2
XOAI21X1_276 INVX1_300/Y INVX1_303/Y AOI22X1_91/C gnd OAI21X1_276/Y vdd OAI21X1
XNAND2X1_390 BUFX2_113/Y AND2X2_8/A gnd OAI21X1_404/B vdd NAND2X1
XNOR2X1_76 gnd INVX1_194/Y gnd NOR2X1_76/Y vdd NOR2X1
XOAI21X1_240 INVX1_262/Y NAND2X1_240/Y OAI21X1_239/Y gnd OAI21X1_240/Y vdd OAI21X1
XNAND2X1_354 BUFX2_41/Y INVX1_401/Y gnd NAND2X1_354/Y vdd NAND2X1
XFILL_28_3_2 gnd vdd FILL
XINVX1_602 INVX1_602/A gnd INVX1_602/Y vdd INVX1
XNAND3X1_186 BUFX2_10/Y INVX1_624/Y INVX1_625/Y gnd NAND3X1_186/Y vdd NAND3X1
XNAND3X1_5 INVX1_5/A OR2X2_5/A NAND3X1_8/C gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_204 INVX1_217/Y OAI21X1_204/B NOR2X1_83/Y gnd AOI21X1_32/C vdd OAI21X1
XNOR2X1_40 INVX1_77/A INVX1_78/Y gnd NOR2X1_40/Y vdd NOR2X1
XNAND2X1_318 INVX1_352/A NAND2X1_317/Y gnd AOI22X1_105/A vdd NAND2X1
XNOR2X1_237 gnd INVX1_600/Y gnd NOR2X1_237/Y vdd NOR2X1
XINVX1_566 INVX1_566/A gnd INVX1_566/Y vdd INVX1
XNAND3X1_150 BUFX2_130/Y INVX1_498/Y INVX1_499/Y gnd NAND3X1_151/B vdd NAND3X1
XCLKBUF1_28 BUFX2_6/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XOAI21X1_168 INVX1_179/Y AOI22X1_54/Y AOI22X1_55/Y gnd OAI21X1_168/Y vdd OAI21X1
XFILL_16_1 gnd vdd FILL
XNOR2X1_201 gnd INVX1_516/Y gnd NOR2X1_201/Y vdd NOR2X1
XNAND2X1_282 INVX1_308/A BUFX2_70/Y gnd NAND2X1_283/B vdd NAND2X1
XNAND3X1_114 BUFX2_118/Y INVX1_372/Y INVX1_373/Y gnd NAND3X1_115/B vdd NAND3X1
XBUFX2_115 NOR3X1_4/Y gnd INVX1_440/A vdd BUFX2
XINVX1_530 BUFX2_33/Y gnd INVX1_530/Y vdd INVX1
XDFFPOSX1_348 INVX1_590/A CLKBUF1_2/Y AOI21X1_85/Y gnd vdd DFFPOSX1
XOAI21X1_132 BUFX2_46/Y INVX1_141/Y INVX1_140/Y gnd OAI21X1_132/Y vdd OAI21X1
XXNOR2X1_75 INVX1_554/A BUFX2_94/Y gnd AOI21X1_80/B vdd XNOR2X1
XNOR2X1_165 gnd INVX1_432/Y gnd NOR2X1_165/Y vdd NOR2X1
XNAND2X1_246 BUFX2_68/Y INVX1_265/Y gnd NAND2X1_246/Y vdd NAND2X1
XDFFPOSX1_312 AND2X2_13/A CLKBUF1_21/Y AOI21X1_76/Y gnd vdd DFFPOSX1
XINVX1_494 INVX1_241/A gnd INVX1_494/Y vdd INVX1
XNOR2X1_129 gnd INVX1_348/Y gnd NOR2X1_129/Y vdd NOR2X1
XXNOR2X1_39 INVX1_293/A BUFX2_52/Y gnd XNOR2X1_39/Y vdd XNOR2X1
XNAND2X1_210 INVX1_219/A NAND2X1_210/B gnd AOI22X1_67/A vdd NAND2X1
XDFFPOSX1_276 INVX1_464/A CLKBUF1_42/Y AOI21X1_67/Y gnd vdd DFFPOSX1
XINVX1_458 INVX1_458/A gnd INVX1_458/Y vdd INVX1
XNAND2X1_174 BUFX2_54/Y INVX1_177/Y gnd AOI22X1_54/D vdd NAND2X1
XDFFPOSX1_240 AND2X2_4/A CLKBUF1_39/Y AOI21X1_58/Y gnd vdd DFFPOSX1
XINVX1_422 INVX1_422/A gnd INVX1_422/Y vdd INVX1
XAOI21X1_72 INVX1_499/Y AOI21X1_72/B AOI21X1_72/C gnd AOI21X1_72/Y vdd AOI21X1
XBUFX2_75 BUFX2_73/A gnd BUFX2_75/Y vdd BUFX2
XNAND2X1_138 BUFX2_50/Y AND2X2_43/B gnd NAND2X1_138/Y vdd NAND2X1
XAOI21X1_36 INVX1_247/Y XNOR2X1_31/Y AOI21X1_36/C gnd AOI21X1_36/Y vdd AOI21X1
XDFFPOSX1_204 INVX1_338/A CLKBUF1_14/Y AOI21X1_49/Y gnd vdd DFFPOSX1
XINVX1_386 BUFX2_37/Y gnd INVX1_386/Y vdd INVX1
XBUFX2_39 BUFX2_39/A gnd BUFX2_39/Y vdd BUFX2
XNAND2X1_99 INVX1_83/A INVX1_86/A gnd OAI21X1_86/B vdd NAND2X1
XOAI21X1_84 BUFX2_76/Y INVX1_83/Y OAI21X1_83/Y gnd OAI21X1_84/Y vdd OAI21X1
XNAND2X1_102 INVX1_84/A BUFX2_76/Y gnd NAND2X1_102/Y vdd NAND2X1
XINVX1_350 NAND2X1_7/A gnd INVX1_350/Y vdd INVX1
XFILL_10_2_0 gnd vdd FILL
XDFFPOSX1_168 INVX1_275/A CLKBUF1_46/Y AOI21X1_40/Y gnd vdd DFFPOSX1
XAOI22X1_170 INVX1_581/A INVX1_580/Y INVX1_582/Y AOI22X1_170/D gnd AOI22X1_170/Y vdd
+ AOI22X1
XOAI21X1_529 INVX1_594/Y INVX1_597/Y AOI22X1_175/C gnd OAI21X1_530/C vdd OAI21X1
XAOI22X1_77 AOI22X1_77/A AND2X2_65/Y AOI22X1_77/C NOR2X1_95/Y gnd AOI22X1_77/Y vdd
+ AOI22X1
XDFFPOSX1_66 AOI22X1_33/C CLKBUF1_1/Y OAI21X1_98/Y gnd vdd DFFPOSX1
XOAI21X1_48 INVX1_41/Y INVX1_44/Y AOI22X1_17/C gnd OAI21X1_48/Y vdd OAI21X1
XDFFPOSX1_132 NAND2X1_9/B CLKBUF1_44/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XNAND2X1_63 INVX1_72/A INVX1_65/A gnd NOR2X1_28/A vdd NAND2X1
XAOI22X1_134 INVX1_455/A INVX1_454/Y INVX1_456/Y NAND2X1_397/Y gnd AOI22X1_134/Y vdd
+ AOI22X1
XOAI21X1_493 INVX1_552/Y INVX1_555/Y OAI21X1_493/C gnd OAI21X1_493/Y vdd OAI21X1
XFILL_16_1_2 gnd vdd FILL
XINVX1_314 INVX1_498/A gnd INVX1_314/Y vdd INVX1
XAOI22X1_41 AOI22X1_41/A AND2X2_44/Y AOI22X1_41/C NOR2X1_56/Y gnd AOI22X1_41/Y vdd
+ AOI22X1
XOAI21X1_12 INVX1_21/Y NOR2X1_17/Y NAND2X1_31/Y gnd OAI21X1_12/Y vdd OAI21X1
XNAND2X1_27 INVX1_5/Y NAND3X1_8/C gnd NAND3X1_12/C vdd NAND2X1
XDFFPOSX1_30 BUFX2_140/A CLKBUF1_28/Y NAND2X1_56/Y gnd vdd DFFPOSX1
XINVX1_278 BUFX2_32/Y gnd INVX1_278/Y vdd INVX1
XAOI21X1_6 XNOR2X1_1/Y XOR2X1_1/Y AOI21X1_6/C gnd AOI21X1_6/Y vdd AOI21X1
XOAI21X1_457 INVX1_510/Y INVX1_513/Y AOI22X1_151/C gnd OAI21X1_458/C vdd OAI21X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XOAI21X1_421 INVX1_468/Y INVX1_471/Y AOI22X1_139/C gnd OAI21X1_421/Y vdd OAI21X1
XNAND3X1_68 INVX1_209/A INVX1_211/Y INVX1_212/Y gnd NAND3X1_69/B vdd NAND3X1
XFILL_17_2_0 gnd vdd FILL
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_206 INVX1_487/A gnd INVX1_206/Y vdd INVX1
XOAI21X1_385 INVX1_426/Y INVX1_429/Y OAI21X1_385/C gnd OAI21X1_386/C vdd OAI21X1
XAND2X2_137 INVX1_601/A INVX1_479/A gnd AND2X2_137/Y vdd AND2X2
XNAND2X1_499 INVX1_597/A INVX1_590/A gnd NOR3X1_8/A vdd NAND2X1
XNAND3X1_32 INVX1_83/A INVX1_85/Y INVX1_86/Y gnd NAND3X1_33/B vdd NAND3X1
XFILL_3_2_2 gnd vdd FILL
XFILL_5_0_1 gnd vdd FILL
XFILL_23_1_2 gnd vdd FILL
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XOAI21X1_349 INVX1_384/Y INVX1_387/Y OAI21X1_349/C gnd OAI21X1_350/C vdd OAI21X1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XAND2X2_101 BUFX2_97/Y INVX1_437/A gnd AND2X2_101/Y vdd AND2X2
XNAND2X1_463 BUFX2_64/Y INVX1_541/Y gnd NAND2X1_463/Y vdd NAND2X1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XAND2X2_74 BUFX2_21/Y AND2X2_74/B gnd AND2X2_74/Y vdd AND2X2
XOAI21X1_313 INVX1_342/Y INVX1_345/Y OAI21X1_313/C gnd OAI21X1_313/Y vdd OAI21X1
XINVX1_134 INVX1_125/A gnd NOR2X1_58/B vdd INVX1
XNAND2X1_427 AND2X2_11/A NAND2X1_427/B gnd AOI22X1_145/A vdd NAND2X1
XAND2X2_38 BUFX2_53/Y INVX1_94/A gnd AND2X2_38/Y vdd AND2X2
XFILL_24_2_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XOAI21X1_277 INVX1_304/Y NAND2X1_274/Y OAI21X1_276/Y gnd OAI21X1_277/Y vdd OAI21X1
XNAND2X1_391 AND2X2_8/Y INVX1_447/Y gnd NAND2X1_391/Y vdd NAND2X1
XNOR2X1_77 AND2X2_8/B NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XOAI21X1_241 INVX1_259/Y OAI21X1_241/B NOR2X1_96/Y gnd AOI21X1_38/C vdd OAI21X1
XNAND2X1_355 INVX1_399/A AND2X2_4/Y gnd NAND2X1_355/Y vdd NAND2X1
XNOR2X1_41 NOR2X1_41/A NOR2X1_41/B gnd BUFX2_103/A vdd NOR2X1
XINVX1_603 BUFX2_11/Y gnd INVX1_603/Y vdd INVX1
XNAND3X1_187 NOR2X1_243/Y NAND3X1_186/Y OAI21X1_552/Y gnd NAND3X1_187/Y vdd NAND3X1
XNAND3X1_6 INVX1_5/A AOI22X1_9/C NAND3X1_8/C gnd NAND3X1_6/Y vdd NAND3X1
XNOR2X1_238 INVX1_602/A INVX1_603/Y gnd NOR2X1_238/Y vdd NOR2X1
XOAI21X1_205 INVX1_221/Y AOI22X1_66/Y AOI22X1_67/Y gnd OAI21X1_205/Y vdd OAI21X1
XNAND2X1_319 BUFX2_122/Y AND2X2_1/A gnd OAI21X1_326/B vdd NAND2X1
XINVX1_567 INVX1_567/A gnd INVX1_567/Y vdd INVX1
XNAND3X1_151 NOR2X1_189/Y NAND3X1_151/B NAND3X1_151/C gnd NAND3X1_151/Y vdd NAND3X1
XCLKBUF1_29 BUFX2_2/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XOAI21X1_169 BUFX2_108/Y NOR2X1_73/B INVX1_182/Y gnd OAI21X1_169/Y vdd OAI21X1
XFILL_16_2 gnd vdd FILL
XNOR2X1_202 INVX1_518/A INVX1_519/Y gnd NOR2X1_202/Y vdd NOR2X1
XNAND2X1_283 INVX1_310/A NAND2X1_283/B gnd AOI22X1_93/A vdd NAND2X1
XDFFPOSX1_349 INVX1_588/A CLKBUF1_2/Y NAND3X1_177/Y gnd vdd DFFPOSX1
XNAND3X1_115 NOR2X1_135/Y NAND3X1_115/B NAND3X1_115/C gnd NAND3X1_115/Y vdd NAND3X1
XBUFX2_116 NOR3X1_4/Y gnd BUFX2_116/Y vdd BUFX2
XINVX1_531 BUFX2_62/Y gnd INVX1_531/Y vdd INVX1
XOAI21X1_133 BUFX2_72/Y INVX1_139/Y OAI21X1_132/Y gnd NAND3X1_49/C vdd OAI21X1
XXNOR2X1_76 BUFX2_125/Y BUFX2_98/Y gnd AOI21X1_81/B vdd XNOR2X1
XNOR2X1_166 INVX1_434/A INVX1_435/Y gnd NOR2X1_166/Y vdd NOR2X1
XNAND2X1_247 BUFX2_60/Y INVX1_268/Y gnd AOI22X1_80/D vdd NAND2X1
XINVX1_495 BUFX2_28/Y gnd INVX1_495/Y vdd INVX1
XDFFPOSX1_313 INVX1_525/A CLKBUF1_26/Y NAND3X1_159/Y gnd vdd DFFPOSX1
XNOR2X1_130 NAND2X1_7/A INVX1_351/Y gnd NOR2X1_130/Y vdd NOR2X1
XXNOR2X1_40 BUFX2_70/Y BUFX2_21/Y gnd AOI21X1_45/B vdd XNOR2X1
XNAND2X1_211 BUFX2_16/Y INVX1_226/A gnd NAND2X1_211/Y vdd NAND2X1
XDFFPOSX1_277 NAND2X1_8/A CLKBUF1_33/Y NAND3X1_141/Y gnd vdd DFFPOSX1
XINVX1_459 INVX1_459/A gnd INVX1_459/Y vdd INVX1
XNAND2X1_175 NOR2X1_71/A INVX1_167/A gnd NAND2X1_175/Y vdd NAND2X1
XDFFPOSX1_241 INVX1_399/A CLKBUF1_39/Y NAND3X1_123/Y gnd vdd DFFPOSX1
XAOI21X1_73 INVX1_506/Y XNOR2X1_68/Y AOI21X1_73/C gnd AOI21X1_73/Y vdd AOI21X1
XINVX1_423 AND2X2_99/B gnd INVX1_423/Y vdd INVX1
XBUFX2_76 BUFX2_73/A gnd BUFX2_76/Y vdd BUFX2
XNAND2X1_139 INVX1_125/A INVX1_132/Y gnd NAND2X1_139/Y vdd NAND2X1
XINVX1_387 INVX1_387/A gnd INVX1_387/Y vdd INVX1
XAOI21X1_37 INVX1_254/Y AOI21X1_37/B AOI21X1_37/C gnd AOI21X1_37/Y vdd AOI21X1
XDFFPOSX1_205 INVX1_336/A CLKBUF1_2/Y NAND3X1_105/Y gnd vdd DFFPOSX1
XBUFX2_40 BUFX2_39/A gnd BUFX2_40/Y vdd BUFX2
XFILL_10_2_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XOAI21X1_85 INVX1_83/Y INVX1_86/Y OAI21X1_85/C gnd OAI21X1_85/Y vdd OAI21X1
XNAND2X1_103 INVX1_86/A NAND2X1_102/Y gnd AOI22X1_29/A vdd NAND2X1
XINVX1_351 BUFX2_118/Y gnd INVX1_351/Y vdd INVX1
XOAI21X1_530 INVX1_598/Y NAND2X1_507/Y OAI21X1_530/C gnd OAI21X1_530/Y vdd OAI21X1
XDFFPOSX1_169 AND2X2_9/B CLKBUF1_20/Y NAND3X1_87/Y gnd vdd DFFPOSX1
XAOI22X1_171 AOI22X1_171/A AND2X2_131/Y OAI21X1_517/C NOR2X1_226/Y gnd AOI22X1_171/Y
+ vdd AOI22X1
XNAND2X1_64 INVX1_56/A INVX1_79/A gnd NOR2X1_28/B vdd NAND2X1
XAOI22X1_78 NOR2X1_97/A INVX1_258/Y INVX1_260/Y AOI22X1_78/D gnd AOI22X1_78/Y vdd
+ AOI22X1
XAOI22X1_135 AOI22X1_135/A AND2X2_104/Y OAI21X1_409/C NOR2X1_172/Y gnd AOI22X1_135/Y
+ vdd AOI22X1
XDFFPOSX1_67 AOI22X1_9/C CLKBUF1_19/Y OAI21X1_100/Y gnd vdd DFFPOSX1
XOAI21X1_49 INVX1_45/Y OAI21X1_49/B OAI21X1_48/Y gnd OAI21X1_49/Y vdd OAI21X1
XDFFPOSX1_133 INVX1_210/A CLKBUF1_5/Y NAND3X1_69/Y gnd vdd DFFPOSX1
XOAI21X1_494 INVX1_556/Y OAI21X1_494/B OAI21X1_493/Y gnd OAI21X1_494/Y vdd OAI21X1
XINVX1_315 AND2X2_12/B gnd INVX1_315/Y vdd INVX1
XAOI22X1_42 INVX1_133/A INVX1_132/Y NOR2X1_58/B AOI22X1_42/D gnd AOI22X1_42/Y vdd
+ AOI22X1
XDFFPOSX1_31 BUFX2_141/A CLKBUF1_6/Y NAND2X1_57/Y gnd vdd DFFPOSX1
XNAND2X1_28 EN_request_put INVX1_17/Y gnd OR2X2_1/A vdd NAND2X1
XOAI21X1_13 INVX1_22/Y NOR2X1_17/Y NAND2X1_32/Y gnd DFFPOSX1_7/D vdd OAI21X1
XAOI21X1_7 INVX1_44/Y AOI21X1_7/B AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_458 INVX1_514/Y OAI21X1_458/B OAI21X1_458/C gnd OAI21X1_458/Y vdd OAI21X1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XINVX1_243 BUFX2_34/Y gnd INVX1_243/Y vdd INVX1
XOAI21X1_422 INVX1_472/Y NAND2X1_408/Y OAI21X1_421/Y gnd OAI21X1_422/Y vdd OAI21X1
XFILL_19_0_0 gnd vdd FILL
XNAND3X1_69 NOR2X1_81/Y NAND3X1_69/B NAND3X1_69/C gnd NAND3X1_69/Y vdd NAND3X1
XFILL_17_2_1 gnd vdd FILL
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XOAI21X1_386 INVX1_430/Y OAI21X1_386/B OAI21X1_386/C gnd OAI21X1_386/Y vdd OAI21X1
XAND2X2_138 BUFX2_11/Y INVX1_612/A gnd AND2X2_138/Y vdd AND2X2
XNAND2X1_500 INVX1_609/A INVX1_604/A gnd NOR3X1_8/B vdd NAND2X1
XNAND3X1_33 NOR2X1_42/Y NAND3X1_33/B OAI21X1_84/Y gnd NAND3X1_33/Y vdd NAND3X1
XFILL_5_0_2 gnd vdd FILL
XINVX1_53 INVX1_45/A gnd INVX1_53/Y vdd INVX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XAND2X2_102 BUFX2_116/Y INVX1_444/A gnd AND2X2_102/Y vdd AND2X2
XOAI21X1_350 INVX1_388/Y OAI21X1_350/B OAI21X1_350/C gnd OAI21X1_350/Y vdd OAI21X1
XNAND2X1_464 INVX1_539/A INVX1_279/A gnd NAND2X1_464/Y vdd NAND2X1
XAND2X2_75 INVX1_498/A INVX1_501/A gnd AND2X2_75/Y vdd AND2X2
XINVX1_17 INVX1_3/Y gnd INVX1_17/Y vdd INVX1
XOAI21X1_314 INVX1_346/Y OAI21X1_314/B OAI21X1_313/Y gnd OAI21X1_314/Y vdd OAI21X1
XINVX1_135 AND2X2_43/B gnd INVX1_135/Y vdd INVX1
XNAND2X1_428 BUFX2_130/Y INVX1_499/A gnd OAI21X1_446/B vdd NAND2X1
XAND2X2_39 BUFX2_105/Y AND2X2_39/B gnd AND2X2_39/Y vdd AND2X2
XFILL_26_0_0 gnd vdd FILL
XNOR3X1_1 INVX1_5/Y NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_4_3_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_24_2_1 gnd vdd FILL
XOAI21X1_278 INVX1_301/Y NAND2X1_275/Y NAND3X1_95/A gnd AOI21X1_44/C vdd OAI21X1
XNAND2X1_392 BUFX2_113/Y INVX1_450/Y gnd AOI22X1_132/D vdd NAND2X1
XNOR2X1_78 gnd NOR2X1_78/B gnd NOR2X1_78/Y vdd NOR2X1
XOAI21X1_242 INVX1_263/Y AOI22X1_78/Y AOI22X1_79/Y gnd OAI21X1_242/Y vdd OAI21X1
XNAND2X1_356 AND2X2_4/A NAND2X1_355/Y gnd NAND2X1_356/Y vdd NAND2X1
XINVX1_604 INVX1_604/A gnd INVX1_604/Y vdd INVX1
XNAND3X1_7 INVX1_5/A OR2X2_3/B NAND3X1_8/C gnd NAND3X1_7/Y vdd NAND3X1
XNOR2X1_42 gnd INVX1_82/Y gnd NOR2X1_42/Y vdd NOR2X1
XOAI21X1_206 BUFX2_15/Y INVX1_225/Y INVX1_224/Y gnd OAI21X1_206/Y vdd OAI21X1
XNOR2X1_239 gnd INVX1_607/Y gnd NOR2X1_239/Y vdd NOR2X1
XNAND2X1_320 AND2X2_1/Y INVX1_356/Y gnd OAI21X1_327/B vdd NAND2X1
XCLKBUF1_30 BUFX2_1/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XINVX1_568 AND2X2_42/A gnd INVX1_568/Y vdd INVX1
XNAND3X1_152 BUFX2_25/Y INVX1_505/Y INVX1_506/Y gnd NAND3X1_152/Y vdd NAND3X1
XOAI21X1_170 BUFX2_67/Y INVX1_181/Y OAI21X1_169/Y gnd NAND3X1_61/C vdd OAI21X1
XNOR2X1_203 gnd INVX1_523/Y gnd NOR2X1_203/Y vdd NOR2X1
XNAND2X1_284 INVX1_319/A INVX1_333/A gnd NAND2X1_284/Y vdd NAND2X1
XDFFPOSX1_350 AOI22X1_175/C CLKBUF1_14/Y OAI21X1_530/Y gnd vdd DFFPOSX1
XNAND3X1_116 BUFX2_75/Y INVX1_379/Y INVX1_380/Y gnd NAND3X1_116/Y vdd NAND3X1
XINVX1_532 INVX1_532/A gnd INVX1_532/Y vdd INVX1
XBUFX2_117 NOR3X1_2/Y gnd BUFX2_117/Y vdd BUFX2
XNOR2X1_167 gnd INVX1_439/Y gnd NOR2X1_167/Y vdd NOR2X1
XOAI21X1_134 INVX1_139/Y INVX1_142/Y AOI22X1_45/C gnd OAI21X1_134/Y vdd OAI21X1
XXNOR2X1_77 AND2X2_42/A INVX1_566/A gnd XNOR2X1_77/Y vdd XNOR2X1
XNAND2X1_248 NOR2X1_99/A BUFX2_68/Y gnd NAND2X1_249/B vdd NAND2X1
XINVX1_496 BUFX2_130/Y gnd INVX1_496/Y vdd INVX1
XDFFPOSX1_314 OAI21X1_475/C CLKBUF1_25/Y OAI21X1_476/Y gnd vdd DFFPOSX1
XXNOR2X1_41 BUFX2_19/Y INVX1_498/A gnd XNOR2X1_41/Y vdd XNOR2X1
XNAND2X1_212 BUFX2_67/Y INVX1_223/Y gnd OAI21X1_210/B vdd NAND2X1
XNOR2X1_131 gnd INVX1_355/Y gnd NOR2X1_131/Y vdd NOR2X1
XDFFPOSX1_278 AOI22X1_139/C CLKBUF1_5/Y OAI21X1_422/Y gnd vdd DFFPOSX1
XINVX1_460 BUFX2_28/Y gnd INVX1_460/Y vdd INVX1
XNAND2X1_176 AND2X2_50/B NAND2X1_175/Y gnd AOI22X1_55/A vdd NAND2X1
XDFFPOSX1_242 AOI22X1_121/C CLKBUF1_27/Y OAI21X1_368/Y gnd vdd DFFPOSX1
XAOI21X1_74 INVX1_513/Y XNOR2X1_69/Y AOI21X1_74/C gnd AOI21X1_74/Y vdd AOI21X1
XINVX1_424 AND2X2_98/B gnd INVX1_424/Y vdd INVX1
XBUFX2_77 BUFX2_73/A gnd BUFX2_77/Y vdd BUFX2
XNAND2X1_140 BUFX2_50/Y INVX1_135/Y gnd AOI22X1_42/D vdd NAND2X1
XINVX1_388 AND2X2_99/B gnd INVX1_388/Y vdd INVX1
XDFFPOSX1_206 OAI21X1_313/C CLKBUF1_41/Y OAI21X1_314/Y gnd vdd DFFPOSX1
XAOI21X1_38 INVX1_261/Y AOI21X1_38/B AOI21X1_38/C gnd AOI21X1_38/Y vdd AOI21X1
XBUFX2_41 BUFX2_39/A gnd BUFX2_41/Y vdd BUFX2
XNAND2X1_104 BUFX2_53/Y INVX1_93/A gnd OAI21X1_92/B vdd NAND2X1
XFILL_10_2_2 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XDFFPOSX1_170 AOI22X1_85/C CLKBUF1_38/Y OAI21X1_259/Y gnd vdd DFFPOSX1
XOAI21X1_86 INVX1_87/Y OAI21X1_86/B OAI21X1_85/Y gnd OAI21X1_86/Y vdd OAI21X1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XAOI22X1_172 INVX1_588/A INVX1_587/Y INVX1_589/Y AOI22X1_172/D gnd OAI21X1_526/B vdd
+ AOI22X1
XOAI21X1_531 INVX1_595/Y NAND2X1_508/Y NOR2X1_235/Y gnd AOI21X1_86/C vdd OAI21X1
XOAI21X1_50 INVX1_42/Y NAND2X1_66/Y NOR2X1_29/Y gnd AOI21X1_7/C vdd OAI21X1
XNAND2X1_65 INVX1_41/A INVX1_44/A gnd OAI21X1_49/B vdd NAND2X1
XAOI22X1_79 AOI22X1_79/A AND2X2_66/Y AOI22X1_79/C NOR2X1_97/Y gnd AOI22X1_79/Y vdd
+ AOI22X1
XAOI22X1_136 NAND2X1_8/A INVX1_461/Y INVX1_463/Y AOI22X1_136/D gnd AOI22X1_136/Y vdd
+ AOI22X1
XDFFPOSX1_68 INVX1_100/A CLKBUF1_19/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 AOI22X1_67/C CLKBUF1_34/Y OAI21X1_203/Y gnd vdd DFFPOSX1
XINVX1_316 BUFX2_18/Y gnd INVX1_316/Y vdd INVX1
XOAI21X1_495 INVX1_553/Y NAND2X1_475/Y NOR2X1_217/Y gnd AOI21X1_80/C vdd OAI21X1
XAOI22X1_43 AOI22X1_43/A AND2X2_45/Y AOI22X1_43/C NOR2X1_58/Y gnd AOI22X1_43/Y vdd
+ AOI22X1
XDFFPOSX1_32 BUFX2_142/A CLKBUF1_28/Y NAND2X1_58/Y gnd vdd DFFPOSX1
XOAI21X1_14 INVX1_23/Y NOR2X1_17/Y NAND2X1_33/Y gnd OAI21X1_14/Y vdd OAI21X1
XNAND2X1_29 request_put[0] NOR2X1_17/Y gnd NAND2X1_29/Y vdd NAND2X1
XFILL_11_3_0 gnd vdd FILL
XOAI21X1_459 INVX1_511/Y OAI21X1_459/B NOR2X1_199/Y gnd AOI21X1_74/C vdd OAI21X1
XAOI21X1_8 INVX1_51/Y XNOR2X1_3/Y AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XAOI22X1_100 INVX1_336/A INVX1_335/Y INVX1_337/Y NAND2X1_306/Y gnd AOI22X1_100/Y vdd
+ AOI22X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XNAND3X1_70 BUFX2_55/Y INVX1_218/Y INVX1_219/Y gnd NAND3X1_71/B vdd NAND3X1
XOAI21X1_423 INVX1_469/Y NAND2X1_409/Y NOR2X1_181/Y gnd AOI21X1_68/C vdd OAI21X1
XFILL_19_0_1 gnd vdd FILL
XFILL_17_2_2 gnd vdd FILL
XOAI21X1_387 INVX1_427/Y OAI21X1_387/B NOR2X1_163/Y gnd AOI21X1_62/C vdd OAI21X1
XINVX1_90 BUFX2_53/Y gnd INVX1_90/Y vdd INVX1
XINVX1_208 BUFX2_30/Y gnd INVX1_208/Y vdd INVX1
XAND2X2_139 BUFX2_13/Y INVX1_619/A gnd AND2X2_139/Y vdd AND2X2
XNAND3X1_34 BUFX2_53/Y INVX1_92/Y INVX1_93/Y gnd NAND3X1_34/Y vdd NAND3X1
XNAND2X1_501 INVX1_623/A INVX1_616/A gnd NOR3X1_8/C vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XINVX1_54 BUFX2_33/Y gnd INVX1_54/Y vdd INVX1
XINVX1_172 INVX1_430/A gnd INVX1_172/Y vdd INVX1
XAND2X2_103 BUFX2_114/Y INVX1_451/A gnd AND2X2_103/Y vdd AND2X2
XOAI21X1_351 INVX1_385/Y OAI21X1_351/B NOR2X1_145/Y gnd AOI21X1_56/C vdd OAI21X1
XNAND2X1_465 AND2X2_15/A NAND2X1_464/Y gnd NAND2X1_465/Y vdd NAND2X1
XAND2X2_76 INVX1_582/A INVX1_325/A gnd AND2X2_76/Y vdd AND2X2
XFILL_18_3_0 gnd vdd FILL
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_429 INVX1_498/A INVX1_496/Y gnd NAND2X1_429/Y vdd NAND2X1
XOAI21X1_315 INVX1_343/Y OAI21X1_315/B NOR2X1_127/Y gnd AOI21X1_50/C vdd OAI21X1
XINVX1_136 OAI21X1_3/Y gnd INVX1_136/Y vdd INVX1
XAND2X2_40 AND2X2_2/Y INVX1_368/A gnd AND2X2_40/Y vdd AND2X2
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XFILL_26_0_1 gnd vdd FILL
XFILL_24_2_2 gnd vdd FILL
XFILL_4_3_2 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XOAI21X1_279 INVX1_305/Y AOI22X1_90/Y AOI22X1_91/Y gnd OAI21X1_279/Y vdd OAI21X1
XNAND2X1_393 INVX1_448/A AND2X2_8/Y gnd NAND2X1_394/B vdd NAND2X1
XNOR2X1_79 AND2X2_10/B NOR2X1_79/B gnd NOR2X1_79/Y vdd NOR2X1
XOAI21X1_243 BUFX2_60/Y NOR2X1_99/B INVX1_266/Y gnd OAI21X1_243/Y vdd OAI21X1
XNAND2X1_357 BUFX2_39/Y AND2X2_5/A gnd OAI21X1_368/B vdd NAND2X1
XINVX1_605 INVX1_479/A gnd INVX1_605/Y vdd INVX1
XOAI21X1_207 BUFX2_69/Y INVX1_223/Y OAI21X1_206/Y gnd NAND3X1_73/C vdd OAI21X1
XNAND3X1_8 INVX1_5/A OR2X2_4/A NAND3X1_8/C gnd OAI21X1_4/C vdd NAND3X1
XNOR2X1_43 INVX1_84/A INVX1_85/Y gnd NOR2X1_43/Y vdd NOR2X1
XFILL_25_3_0 gnd vdd FILL
XNOR2X1_240 INVX1_609/A INVX1_610/Y gnd NOR2X1_240/Y vdd NOR2X1
XNAND2X1_321 BUFX2_122/Y INVX1_359/Y gnd NAND2X1_321/Y vdd NAND2X1
XCLKBUF1_31 BUFX2_5/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XINVX1_569 AND2X2_16/A gnd INVX1_569/Y vdd INVX1
XNAND3X1_153 NOR2X1_197/Y NAND3X1_152/Y NAND3X1_153/C gnd NAND3X1_153/Y vdd NAND3X1
XOAI21X1_171 INVX1_181/Y INVX1_184/Y AOI22X1_57/C gnd OAI21X1_172/C vdd OAI21X1
XNOR2X1_204 INVX1_525/A INVX1_526/Y gnd NOR2X1_204/Y vdd NOR2X1
XNAND2X1_285 NAND2X1_284/Y OAI21X1_286/Y gnd AND2X2_74/B vdd NAND2X1
XNAND3X1_117 NOR2X1_143/Y NAND3X1_116/Y OAI21X1_342/Y gnd NAND3X1_117/Y vdd NAND3X1
XINVX1_533 INVX1_244/A gnd INVX1_533/Y vdd INVX1
XDFFPOSX1_351 INVX1_599/A CLKBUF1_14/Y OAI21X1_532/Y gnd vdd DFFPOSX1
XBUFX2_118 NOR3X1_2/Y gnd BUFX2_118/Y vdd BUFX2
XNOR2X1_168 INVX1_441/A INVX1_442/Y gnd NOR2X1_168/Y vdd NOR2X1
XOAI21X1_135 INVX1_143/Y NAND2X1_143/Y OAI21X1_134/Y gnd OAI21X1_135/Y vdd OAI21X1
XXNOR2X1_78 INVX1_575/A BUFX2_124/Y gnd XNOR2X1_78/Y vdd XNOR2X1
XNAND2X1_249 INVX1_268/A NAND2X1_249/B gnd AOI22X1_81/A vdd NAND2X1
XINVX1_497 INVX1_497/A gnd INVX1_497/Y vdd INVX1
XDFFPOSX1_315 AND2X2_63/B CLKBUF1_29/Y OAI21X1_478/Y gnd vdd DFFPOSX1
XXNOR2X1_42 BUFX2_18/Y INVX1_582/A gnd XNOR2X1_42/Y vdd XNOR2X1
XNAND2X1_213 BUFX2_15/Y INVX1_226/Y gnd AOI22X1_68/D vdd NAND2X1
XNOR2X1_132 INVX1_357/A INVX1_358/Y gnd NOR2X1_132/Y vdd NOR2X1
XDFFPOSX1_279 INVX1_473/A CLKBUF1_25/Y OAI21X1_424/Y gnd vdd DFFPOSX1
XINVX1_461 BUFX2_83/Y gnd INVX1_461/Y vdd INVX1
XNAND2X1_177 BUFX2_108/Y INVX1_184/A gnd OAI21X1_172/B vdd NAND2X1
XDFFPOSX1_243 AND2X2_47/B CLKBUF1_27/Y OAI21X1_370/Y gnd vdd DFFPOSX1
XINVX1_425 BUFX2_34/Y gnd INVX1_425/Y vdd INVX1
XAOI21X1_75 INVX1_520/Y XNOR2X1_70/Y AOI21X1_75/C gnd AOI21X1_75/Y vdd AOI21X1
XBUFX2_78 BUFX2_79/A gnd BUFX2_78/Y vdd BUFX2
XNAND2X1_141 INVX1_133/A INVX1_125/A gnd NAND2X1_141/Y vdd NAND2X1
XDFFPOSX1_207 AND2X2_80/A CLKBUF1_48/Y OAI21X1_316/Y gnd vdd DFFPOSX1
XINVX1_389 AND2X2_87/B gnd INVX1_389/Y vdd INVX1
XAOI21X1_39 INVX1_268/Y AOI21X1_39/B AOI21X1_39/C gnd AOI21X1_39/Y vdd AOI21X1
XFILL_20_1 gnd vdd FILL
XBUFX2_42 BUFX2_44/A gnd BUFX2_42/Y vdd BUFX2
XFILL_12_0_2 gnd vdd FILL
XNAND2X1_105 INVX1_83/A INVX1_90/Y gnd OAI21X1_93/B vdd NAND2X1
XDFFPOSX1_171 INVX1_284/A CLKBUF1_46/Y OAI21X1_261/Y gnd vdd DFFPOSX1
XAOI22X1_173 AOI22X1_173/A AND2X2_135/Y AOI22X1_173/C NOR2X1_234/Y gnd OAI21X1_526/C
+ vdd AOI22X1
XOAI21X1_87 INVX1_84/Y OAI21X1_87/B NOR2X1_42/Y gnd OAI21X1_87/Y vdd OAI21X1
XINVX1_353 INVX1_430/A gnd INVX1_353/Y vdd INVX1
XOAI21X1_532 INVX1_599/Y AOI22X1_174/Y AOI22X1_175/Y gnd OAI21X1_532/Y vdd OAI21X1
XAOI22X1_80 NOR2X1_99/A INVX1_265/Y NOR2X1_99/B AOI22X1_80/D gnd AOI22X1_80/Y vdd
+ AOI22X1
XDFFPOSX1_69 INVX1_98/A CLKBUF1_19/Y NAND3X1_37/Y gnd vdd DFFPOSX1
XNAND2X1_66 INVX1_43/A INVX1_41/Y gnd NAND2X1_66/Y vdd NAND2X1
XOAI21X1_51 INVX1_46/Y OAI21X1_51/B OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XAOI22X1_137 AOI22X1_137/A AND2X2_108/Y AOI22X1_137/C NOR2X1_180/Y gnd AOI22X1_137/Y
+ vdd AOI22X1
XOAI21X1_496 INVX1_557/Y OAI21X1_496/B OAI21X1_496/C gnd OAI21X1_496/Y vdd OAI21X1
XDFFPOSX1_135 INVX1_221/A CLKBUF1_34/Y OAI21X1_205/Y gnd vdd DFFPOSX1
XINVX1_317 INVX1_317/A gnd INVX1_317/Y vdd INVX1
XAOI22X1_44 INVX1_140/A INVX1_139/Y INVX1_141/Y AOI22X1_44/D gnd AOI22X1_44/Y vdd
+ AOI22X1
XDFFPOSX1_33 BUFX2_143/A CLKBUF1_28/Y NAND2X1_59/Y gnd vdd DFFPOSX1
XNAND2X1_30 request_put[1] NOR2X1_17/Y gnd OAI21X1_11/C vdd NAND2X1
XOAI21X1_15 INVX1_24/Y NOR2X1_17/Y OAI21X1_15/C gnd DFFPOSX1_9/D vdd OAI21X1
XFILL_11_3_1 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XOAI21X1_460 INVX1_515/Y OAI21X1_460/B AOI22X1_151/Y gnd OAI21X1_460/Y vdd OAI21X1
XINVX1_281 BUFX2_59/Y gnd INVX1_281/Y vdd INVX1
XAOI21X1_9 INVX1_58/Y AOI21X1_9/B AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XAOI22X1_101 AOI22X1_101/A AND2X2_81/Y OAI21X1_307/C NOR2X1_126/Y gnd OAI21X1_310/C
+ vdd AOI22X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XNAND3X1_71 NOR2X1_83/Y NAND3X1_71/B NAND3X1_71/C gnd NAND3X1_71/Y vdd NAND3X1
XOAI21X1_424 INVX1_473/Y OAI21X1_424/B OAI21X1_424/C gnd OAI21X1_424/Y vdd OAI21X1
XFILL_19_0_2 gnd vdd FILL
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XOAI21X1_388 INVX1_431/Y AOI22X1_126/Y AOI22X1_127/Y gnd OAI21X1_388/Y vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XAND2X2_140 BUFX2_10/Y INVX1_626/A gnd AND2X2_140/Y vdd AND2X2
XNAND3X1_35 NOR2X1_44/Y NAND3X1_34/Y OAI21X1_90/Y gnd NAND3X1_35/Y vdd NAND3X1
XNAND2X1_502 BUFX2_26/Y INVX1_590/A gnd NAND2X1_502/Y vdd NAND2X1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XAND2X2_104 BUFX2_112/Y INVX1_458/A gnd AND2X2_104/Y vdd AND2X2
XOAI21X1_352 INVX1_389/Y OAI21X1_352/B AOI22X1_115/Y gnd OAI21X1_352/Y vdd OAI21X1
XINVX1_173 BUFX2_30/Y gnd NOR2X1_70/B vdd INVX1
XNAND2X1_466 INVX1_555/A INVX1_548/A gnd NOR3X1_7/A vdd NAND2X1
XFILL_20_1_0 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XAND2X2_77 INVX1_624/A INVX1_627/A gnd AND2X2_77/Y vdd AND2X2
XFILL_18_3_1 gnd vdd FILL
XOAI21X1_316 INVX1_347/Y OAI21X1_316/B AOI22X1_103/Y gnd OAI21X1_316/Y vdd OAI21X1
XINVX1_19 OR2X2_1/B gnd INVX1_19/Y vdd INVX1
XINVX1_137 INVX1_129/A gnd INVX1_137/Y vdd INVX1
XNAND2X1_430 BUFX2_130/Y INVX1_499/Y gnd AOI22X1_146/D vdd NAND2X1
XAND2X2_41 AND2X2_4/Y INVX1_115/A gnd AND2X2_41/Y vdd AND2X2
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd BUFX2_39/A vdd NOR3X1
XFILL_6_1_2 gnd vdd FILL
XFILL_26_0_2 gnd vdd FILL
XINVX1_101 AND2X2_39/B gnd INVX1_101/Y vdd INVX1
XOAI21X1_280 BUFX2_21/Y INVX1_309/Y INVX1_308/Y gnd OAI21X1_281/C vdd OAI21X1
XNAND2X1_394 AND2X2_8/A NAND2X1_394/B gnd AOI22X1_133/A vdd NAND2X1
XNOR2X1_80 NOR2X1_80/A NOR2X1_80/B gnd BUFX2_17/A vdd NOR2X1
XOAI21X1_244 BUFX2_68/Y INVX1_265/Y OAI21X1_243/Y gnd NAND3X1_85/C vdd OAI21X1
XNAND2X1_358 AND2X2_5/Y INVX1_405/Y gnd NAND2X1_358/Y vdd NAND2X1
XINVX1_606 INVX1_606/A gnd INVX1_606/Y vdd INVX1
XNAND3X1_9 INVX1_5/A OR2X2_4/B NAND3X1_8/C gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_208 INVX1_223/Y INVX1_226/Y AOI22X1_69/C gnd OAI21X1_209/C vdd OAI21X1
XNOR2X1_44 gnd INVX1_89/Y gnd NOR2X1_44/Y vdd NOR2X1
XFILL_27_1_0 gnd vdd FILL
XFILL_25_3_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XNOR2X1_241 gnd INVX1_614/Y gnd NOR2X1_241/Y vdd NOR2X1
XNAND2X1_322 INVX1_357/A AND2X2_1/Y gnd NAND2X1_323/B vdd NAND2X1
XINVX1_570 INVX1_570/A gnd INVX1_570/Y vdd INVX1
XCLKBUF1_32 BUFX2_2/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XNAND3X1_154 BUFX2_89/Y INVX1_512/Y INVX1_513/Y gnd NAND3X1_154/Y vdd NAND3X1
XOAI21X1_172 INVX1_185/Y OAI21X1_172/B OAI21X1_172/C gnd OAI21X1_172/Y vdd OAI21X1
XNOR2X1_205 gnd INVX1_530/Y gnd NOR2X1_205/Y vdd NOR2X1
XNAND2X1_286 INVX1_498/A INVX1_317/A gnd OAI21X1_290/B vdd NAND2X1
XBUFX2_119 NOR3X1_2/Y gnd INVX1_363/A vdd BUFX2
XNAND3X1_118 BUFX2_79/Y INVX1_386/Y INVX1_387/Y gnd NAND3X1_119/B vdd NAND3X1
XDFFPOSX1_352 INVX1_597/A CLKBUF1_50/Y AOI21X1_86/Y gnd vdd DFFPOSX1
XINVX1_534 AND2X2_14/A gnd INVX1_534/Y vdd INVX1
XXNOR2X1_79 INVX1_582/A INVX1_580/A gnd XNOR2X1_79/Y vdd XNOR2X1
XOAI21X1_136 INVX1_140/Y OAI21X1_136/B NOR2X1_59/Y gnd AOI21X1_21/C vdd OAI21X1
XNOR2X1_169 gnd INVX1_446/Y gnd NOR2X1_169/Y vdd NOR2X1
XNAND2X1_250 INVX1_277/A INVX1_291/A gnd NAND2X1_251/A vdd NAND2X1
XDFFPOSX1_316 AND2X2_14/A CLKBUF1_11/Y AOI21X1_77/Y gnd vdd DFFPOSX1
XINVX1_498 INVX1_498/A gnd INVX1_498/Y vdd INVX1
XOAI21X1_100 INVX1_102/Y AOI22X1_32/Y AOI22X1_33/Y gnd OAI21X1_100/Y vdd OAI21X1
XXNOR2X1_43 BUFX2_20/Y INVX1_624/A gnd XNOR2X1_43/Y vdd XNOR2X1
XNOR2X1_133 gnd INVX1_362/Y gnd NOR2X1_133/Y vdd NOR2X1
XNAND2X1_214 INVX1_224/A BUFX2_69/Y gnd NAND2X1_214/Y vdd NAND2X1
XINVX1_462 NAND2X1_8/A gnd INVX1_462/Y vdd INVX1
XDFFPOSX1_280 INVX1_471/A CLKBUF1_25/Y AOI21X1_68/Y gnd vdd DFFPOSX1
XNAND2X1_178 BUFX2_67/Y INVX1_181/Y gnd OAI21X1_173/B vdd NAND2X1
XINVX1_426 BUFX2_84/Y gnd INVX1_426/Y vdd INVX1
XDFFPOSX1_244 AND2X2_5/A CLKBUF1_30/Y AOI21X1_59/Y gnd vdd DFFPOSX1
XAOI21X1_76 INVX1_527/Y AOI21X1_76/B AOI21X1_76/C gnd AOI21X1_76/Y vdd AOI21X1
XBUFX2_79 BUFX2_79/A gnd BUFX2_79/Y vdd BUFX2
XNAND2X1_142 AND2X2_43/B NAND2X1_141/Y gnd AOI22X1_43/A vdd NAND2X1
XDFFPOSX1_208 INVX1_345/A CLKBUF1_41/Y AOI21X1_50/Y gnd vdd DFFPOSX1
XAOI21X1_40 INVX1_275/Y XNOR2X1_35/Y AOI21X1_40/C gnd AOI21X1_40/Y vdd AOI21X1
XINVX1_390 BUFX2_30/Y gnd INVX1_390/Y vdd INVX1
XFILL_20_2 gnd vdd FILL
XBUFX2_43 BUFX2_44/A gnd BUFX2_43/Y vdd BUFX2
XNAND2X1_106 BUFX2_53/Y INVX1_93/Y gnd AOI22X1_30/D vdd NAND2X1
XOAI21X1_88 INVX1_88/Y OAI21X1_88/B OAI21X1_88/C gnd OAI21X1_88/Y vdd OAI21X1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XOAI21X1_533 BUFX2_99/Y INVX1_603/Y INVX1_602/Y gnd OAI21X1_534/C vdd OAI21X1
XDFFPOSX1_172 INVX1_282/A CLKBUF1_46/Y AOI21X1_41/Y gnd vdd DFFPOSX1
XAOI22X1_174 NAND2X1_6/B INVX1_594/Y INVX1_596/Y NAND2X1_509/Y gnd AOI22X1_174/Y vdd
+ AOI22X1
XAOI22X1_81 AOI22X1_81/A AND2X2_67/Y AOI22X1_81/C NOR2X1_99/Y gnd AOI22X1_81/Y vdd
+ AOI22X1
XDFFPOSX1_70 AOI22X1_35/C CLKBUF1_43/Y DFFPOSX1_70/D gnd vdd DFFPOSX1
XNAND2X1_67 INVX1_41/A INVX1_44/Y gnd AOI22X1_16/D vdd NAND2X1
XOAI21X1_52 BUFX2_56/Y INVX1_50/Y INVX1_49/Y gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_497 BUFX2_98/Y INVX1_561/Y INVX1_560/Y gnd OAI21X1_497/Y vdd OAI21X1
XINVX1_318 INVX1_501/A gnd INVX1_318/Y vdd INVX1
XDFFPOSX1_136 INVX1_219/A CLKBUF1_12/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XAOI22X1_138 INVX1_469/A INVX1_468/Y INVX1_470/Y AOI22X1_138/D gnd OAI21X1_424/B vdd
+ AOI22X1
XAOI22X1_45 AOI22X1_45/A AND2X2_46/Y AOI22X1_45/C NOR2X1_60/Y gnd AOI22X1_45/Y vdd
+ AOI22X1
XNAND2X1_31 request_put[2] NOR2X1_17/Y gnd NAND2X1_31/Y vdd NAND2X1
XDFFPOSX1_100 INVX1_156/A CLKBUF1_43/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XFILL_13_1_1 gnd vdd FILL
XAOI22X1_102 INVX1_343/A INVX1_342/Y INVX1_344/Y NAND2X1_311/Y gnd OAI21X1_316/B vdd
+ AOI22X1
XOAI21X1_16 INVX1_25/Y NOR2X1_17/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XDFFPOSX1_34 AOI22X1_17/C CLKBUF1_24/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XFILL_11_3_2 gnd vdd FILL
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XOAI21X1_461 BUFX2_93/Y INVX1_519/Y INVX1_518/Y gnd OAI21X1_461/Y vdd OAI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XINVX1_246 BUFX2_15/Y gnd NOR2X1_92/B vdd INVX1
XOAI21X1_425 INVX1_475/A INVX1_477/Y INVX1_476/Y gnd OAI21X1_425/Y vdd OAI21X1
XNAND3X1_72 BUFX2_16/Y INVX1_225/Y INVX1_226/Y gnd NAND3X1_73/B vdd NAND3X1
XINVX1_92 INVX1_83/A gnd INVX1_92/Y vdd INVX1
XOAI21X1_389 BUFX2_96/Y INVX1_435/Y INVX1_434/Y gnd OAI21X1_389/Y vdd OAI21X1
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XNAND3X1_36 INVX1_97/A INVX1_99/Y INVX1_100/Y gnd NAND3X1_36/Y vdd NAND3X1
XNAND2X1_503 BUFX2_12/Y INVX1_587/Y gnd OAI21X1_525/B vdd NAND2X1
XINVX1_174 BUFX2_54/Y gnd INVX1_174/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XAND2X2_105 INVX1_480/A INVX1_473/A gnd NOR2X1_174/B vdd AND2X2
XNAND2X1_467 INVX1_567/A INVX1_562/A gnd NOR3X1_7/B vdd NAND2X1
XOAI21X1_353 BUFX2_88/Y INVX1_393/Y INVX1_392/Y gnd OAI21X1_354/C vdd OAI21X1
XFILL_2_0_0 gnd vdd FILL
XFILL_20_1_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XAND2X2_78 INVX1_354/A AND2X2_80/A gnd AND2X2_78/Y vdd AND2X2
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XFILL_18_3_2 gnd vdd FILL
XOAI21X1_317 BUFX2_86/Y INVX1_351/Y INVX1_350/Y gnd OAI21X1_317/Y vdd OAI21X1
XINVX1_138 BUFX2_28/Y gnd NOR2X1_59/B vdd INVX1
XNAND2X1_431 INVX1_497/A INVX1_498/A gnd NAND2X1_432/B vdd NAND2X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XAND2X2_42 AND2X2_42/A INVX1_122/A gnd AND2X2_42/Y vdd AND2X2
XINVX1_102 AOI22X1_9/C gnd INVX1_102/Y vdd INVX1
XOAI21X1_281 INVX1_99/A INVX1_307/Y OAI21X1_281/C gnd NAND3X1_97/C vdd OAI21X1
XNAND2X1_395 BUFX2_114/Y AND2X2_9/A gnd OAI21X1_410/B vdd NAND2X1
XNOR2X1_81 gnd INVX1_208/Y gnd NOR2X1_81/Y vdd NOR2X1
XOAI21X1_245 INVX1_265/Y INVX1_268/Y AOI22X1_81/C gnd OAI21X1_246/C vdd OAI21X1
XNAND2X1_359 BUFX2_39/Y INVX1_408/Y gnd NAND2X1_359/Y vdd NAND2X1
XFILL_11_1 gnd vdd FILL
XINVX1_607 BUFX2_30/Y gnd INVX1_607/Y vdd INVX1
XOAI21X1_209 INVX1_227/Y NAND2X1_211/Y OAI21X1_209/C gnd OAI21X1_209/Y vdd OAI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XFILL_27_1_1 gnd vdd FILL
XFILL_25_3_2 gnd vdd FILL
XNOR2X1_45 INVX1_91/A INVX1_92/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_242 INVX1_616/A INVX1_617/Y gnd NOR2X1_242/Y vdd NOR2X1
XNAND2X1_323 AND2X2_1/A NAND2X1_323/B gnd AOI22X1_107/A vdd NAND2X1
XCLKBUF1_33 BUFX2_1/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XINVX1_571 INVX1_122/A gnd INVX1_571/Y vdd INVX1
XNAND3X1_155 NOR2X1_199/Y NAND3X1_154/Y OAI21X1_456/Y gnd NAND3X1_155/Y vdd NAND3X1
XOAI21X1_173 INVX1_182/Y OAI21X1_173/B NOR2X1_72/Y gnd AOI21X1_27/C vdd OAI21X1
XNOR2X1_206 INVX1_532/A INVX1_533/Y gnd NOR2X1_206/Y vdd NOR2X1
XNAND2X1_287 BUFX2_18/Y INVX1_314/Y gnd NAND2X1_287/Y vdd NAND2X1
XBUFX2_120 NOR3X1_2/Y gnd AND2X2_85/A vdd BUFX2
XNAND3X1_119 NOR2X1_145/Y NAND3X1_119/B NAND3X1_119/C gnd NAND3X1_119/Y vdd NAND3X1
XDFFPOSX1_353 NAND2X1_6/B CLKBUF1_50/Y NAND3X1_179/Y gnd vdd DFFPOSX1
XINVX1_535 INVX1_535/A gnd INVX1_535/Y vdd INVX1
XOAI21X1_137 INVX1_144/Y AOI22X1_44/Y AOI22X1_45/Y gnd OAI21X1_137/Y vdd OAI21X1
XXNOR2X1_80 BUFX2_12/Y BUFX2_26/Y gnd AOI21X1_85/B vdd XNOR2X1
XNOR2X1_170 INVX1_448/A INVX1_449/Y gnd NOR2X1_170/Y vdd NOR2X1
XNAND2X1_251 NAND2X1_251/A NAND2X1_251/B gnd INVX1_269/A vdd NAND2X1
XDFFPOSX1_317 INVX1_532/A CLKBUF1_11/Y NAND3X1_161/Y gnd vdd DFFPOSX1
XINVX1_499 INVX1_499/A gnd INVX1_499/Y vdd INVX1
XNOR2X1_134 INVX1_364/A INVX1_365/Y gnd NOR2X1_134/Y vdd NOR2X1
XOAI21X1_101 INVX1_109/A INVX1_123/A INVX1_116/A gnd OAI21X1_101/Y vdd OAI21X1
XXNOR2X1_44 BUFX2_117/Y BUFX2_22/Y gnd AOI21X1_49/B vdd XNOR2X1
XNAND2X1_215 INVX1_226/A NAND2X1_214/Y gnd AOI22X1_69/A vdd NAND2X1
XINVX1_463 INVX1_463/A gnd INVX1_463/Y vdd INVX1
XDFFPOSX1_281 INVX1_469/A CLKBUF1_21/Y NAND3X1_143/Y gnd vdd DFFPOSX1
XNAND2X1_179 BUFX2_108/Y INVX1_184/Y gnd AOI22X1_56/D vdd NAND2X1
XDFFPOSX1_245 INVX1_406/A CLKBUF1_27/Y NAND3X1_125/Y gnd vdd DFFPOSX1
XINVX1_427 INVX1_427/A gnd INVX1_427/Y vdd INVX1
XAOI21X1_77 INVX1_534/Y XNOR2X1_72/Y AOI21X1_77/C gnd AOI21X1_77/Y vdd AOI21X1
XBUFX2_80 BUFX2_79/A gnd BUFX2_80/Y vdd BUFX2
XNAND2X1_143 BUFX2_46/Y INVX1_142/A gnd NAND2X1_143/Y vdd NAND2X1
XAOI21X1_41 INVX1_282/Y AOI21X1_41/B AOI21X1_41/C gnd AOI21X1_41/Y vdd AOI21X1
XDFFPOSX1_209 INVX1_343/A CLKBUF1_48/Y NAND3X1_107/Y gnd vdd DFFPOSX1
XINVX1_391 BUFX2_88/Y gnd INVX1_391/Y vdd INVX1
XBUFX2_44 BUFX2_44/A gnd INVX1_64/A vdd BUFX2
XOAI21X1_89 BUFX2_53/Y INVX1_92/Y INVX1_91/Y gnd OAI21X1_89/Y vdd OAI21X1
XNAND2X1_107 INVX1_91/A INVX1_83/A gnd NAND2X1_108/B vdd NAND2X1
XOAI21X1_534 BUFX2_11/Y INVX1_601/Y OAI21X1_534/C gnd NAND3X1_181/C vdd OAI21X1
XAOI22X1_175 NAND2X1_511/Y AND2X2_136/Y AOI22X1_175/C NOR2X1_236/Y gnd AOI22X1_175/Y
+ vdd AOI22X1
XDFFPOSX1_173 INVX1_280/A CLKBUF1_22/Y NAND3X1_89/Y gnd vdd DFFPOSX1
XINVX1_355 BUFX2_30/Y gnd INVX1_355/Y vdd INVX1
XAOI22X1_82 AND2X2_9/B INVX1_272/Y INVX1_274/Y AOI22X1_82/D gnd AOI22X1_82/Y vdd AOI22X1
XDFFPOSX1_71 INVX1_109/A CLKBUF1_15/Y OAI21X1_107/Y gnd vdd DFFPOSX1
XNAND2X1_68 INVX1_42/A BUFX2_24/Y gnd NAND2X1_68/Y vdd NAND2X1
XOAI21X1_53 INVX1_41/A INVX1_48/Y OAI21X1_52/Y gnd OAI21X1_53/Y vdd OAI21X1
XDFFPOSX1_137 INVX1_217/A CLKBUF1_44/Y NAND3X1_71/Y gnd vdd DFFPOSX1
XOAI21X1_498 BUFX2_125/Y INVX1_559/Y OAI21X1_497/Y gnd NAND3X1_169/C vdd OAI21X1
XAOI22X1_139 NAND2X1_412/Y AND2X2_109/Y AOI22X1_139/C NOR2X1_182/Y gnd OAI21X1_424/C
+ vdd AOI22X1
XINVX1_319 INVX1_319/A gnd INVX1_319/Y vdd INVX1
XAOI22X1_46 AND2X2_5/B INVX1_146/Y NOR2X1_62/B AOI22X1_46/D gnd AOI22X1_46/Y vdd AOI22X1
XOAI21X1_17 INVX1_16/Y AND2X2_23/B NOR2X1_16/Y gnd AOI21X1_1/C vdd OAI21X1
XNAND2X1_32 request_put[3] NOR2X1_17/Y gnd NAND2X1_32/Y vdd NAND2X1
XDFFPOSX1_101 AND2X2_7/B CLKBUF1_43/Y NAND3X1_53/Y gnd vdd DFFPOSX1
XFILL_13_1_2 gnd vdd FILL
XAOI22X1_103 AOI22X1_103/A AND2X2_82/Y OAI21X1_313/C NOR2X1_128/Y gnd AOI22X1_103/Y
+ vdd AOI22X1
XDFFPOSX1_35 INVX1_46/A CLKBUF1_24/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XOAI21X1_462 BUFX2_65/Y INVX1_517/Y OAI21X1_461/Y gnd OAI21X1_462/Y vdd OAI21X1
XAOI22X1_10 INVX1_33/A AOI22X1_9/B OR2X2_3/B AOI22X1_9/D gnd AOI22X1_10/Y vdd AOI22X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XOAI21X1_426 BUFX2_133/Y INVX1_475/Y OAI21X1_425/Y gnd OAI21X1_426/Y vdd OAI21X1
XNAND3X1_73 NOR2X1_85/Y NAND3X1_73/B NAND3X1_73/C gnd NAND3X1_73/Y vdd NAND3X1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XOAI21X1_390 BUFX2_112/Y INVX1_433/Y OAI21X1_389/Y gnd NAND3X1_133/C vdd OAI21X1
XNAND3X1_37 NOR2X1_46/Y NAND3X1_36/Y OAI21X1_96/Y gnd NAND3X1_37/Y vdd NAND3X1
XFILL_14_2_0 gnd vdd FILL
XINVX1_211 BUFX2_91/Y gnd INVX1_211/Y vdd INVX1
XNAND2X1_504 BUFX2_26/Y INVX1_590/Y gnd AOI22X1_172/D vdd NAND2X1
XINVX1_175 NOR2X1_71/A gnd INVX1_175/Y vdd INVX1
XOAI21X1_354 BUFX2_36/Y INVX1_391/Y OAI21X1_354/C gnd NAND3X1_121/C vdd OAI21X1
XINVX1_57 BUFX2_70/Y gnd INVX1_57/Y vdd INVX1
XAND2X2_106 INVX1_480/A INVX1_466/A gnd NOR2X1_176/B vdd AND2X2
XNAND2X1_468 INVX1_581/A INVX1_574/A gnd NOR3X1_7/C vdd NAND2X1
XFILL_2_0_1 gnd vdd FILL
XAND2X2_79 INVX1_354/A AND2X2_79/B gnd AND2X2_79/Y vdd AND2X2
XFILL_20_1_2 gnd vdd FILL
XFILL_0_2_2 gnd vdd FILL
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_139 BUFX2_46/Y gnd INVX1_139/Y vdd INVX1
XOAI21X1_318 BUFX2_118/Y INVX1_349/Y OAI21X1_317/Y gnd NAND3X1_109/C vdd OAI21X1
XNAND2X1_432 INVX1_499/A NAND2X1_432/B gnd AOI22X1_147/A vdd NAND2X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XAND2X2_43 NOR2X1_56/A AND2X2_43/B gnd INVX1_125/A vdd AND2X2
XINVX1_103 BUFX2_35/Y gnd INVX1_103/Y vdd INVX1
XNAND2X1_396 AND2X2_9/Y INVX1_454/Y gnd OAI21X1_411/B vdd NAND2X1
XAOI22X1_1 INVX1_18/A AOI22X1_4/B request_put[0] AOI22X1_4/D gnd AOI22X1_1/Y vdd AOI22X1
XOAI21X1_282 INVX1_307/Y INVX1_310/Y AOI22X1_93/C gnd OAI21X1_283/C vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XNOR2X1_82 INVX1_210/A INVX1_211/Y gnd NOR2X1_82/Y vdd NOR2X1
XOAI21X1_246 INVX1_269/Y NAND2X1_245/Y OAI21X1_246/C gnd OAI21X1_246/Y vdd OAI21X1
XNAND2X1_360 INVX1_406/A AND2X2_5/Y gnd NAND2X1_361/B vdd NAND2X1
XFILL_11_2 gnd vdd FILL
XNOR2X1_46 gnd INVX1_96/Y gnd NOR2X1_46/Y vdd NOR2X1
XFILL_27_1_2 gnd vdd FILL
XINVX1_608 BUFX2_9/Y gnd INVX1_608/Y vdd INVX1
XOAI21X1_210 INVX1_224/Y OAI21X1_210/B NOR2X1_85/Y gnd AOI21X1_33/C vdd OAI21X1
XFILL_7_2_2 gnd vdd FILL
XFILL_9_0_1 gnd vdd FILL
XNOR2X1_243 gnd INVX1_621/Y gnd NOR2X1_243/Y vdd NOR2X1
XNAND2X1_324 INVX1_363/A AND2X2_2/A gnd OAI21X1_332/B vdd NAND2X1
XCLKBUF1_34 BUFX2_7/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XINVX1_572 BUFX2_32/Y gnd INVX1_572/Y vdd INVX1
XNAND3X1_156 BUFX2_93/Y INVX1_519/Y INVX1_520/Y gnd NAND3X1_156/Y vdd NAND3X1
XOAI21X1_174 INVX1_186/Y AOI22X1_56/Y AOI22X1_57/Y gnd OAI21X1_174/Y vdd OAI21X1
XNOR2X1_10 NOR2X1_10/A INVX1_4/Y gnd NAND3X1_3/B vdd NOR2X1
XXNOR2X1_1 AOI22X1_9/C INVX1_39/A gnd XNOR2X1_1/Y vdd XNOR2X1
XNOR2X1_207 gnd INVX1_537/Y gnd NOR2X1_207/Y vdd NOR2X1
XNAND2X1_288 INVX1_498/A INVX1_317/Y gnd AOI22X1_94/D vdd NAND2X1
XDFFPOSX1_354 OAI21X1_535/C CLKBUF1_32/Y OAI21X1_536/Y gnd vdd DFFPOSX1
XBUFX2_121 NOR3X1_2/Y gnd INVX1_370/A vdd BUFX2
XNAND3X1_120 BUFX2_88/Y INVX1_393/Y INVX1_394/Y gnd NAND3X1_121/B vdd NAND3X1
XINVX1_536 AND2X2_63/B gnd INVX1_536/Y vdd INVX1
XOAI21X1_138 INVX1_151/A INVX1_165/A INVX1_158/A gnd OAI21X1_138/Y vdd OAI21X1
XXNOR2X1_81 BUFX2_13/Y BUFX2_78/Y gnd XNOR2X1_81/Y vdd XNOR2X1
XFILL_28_2_0 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XNOR2X1_171 gnd INVX1_453/Y gnd NOR2X1_171/Y vdd NOR2X1
XNAND2X1_252 AND2X2_9/Y INVX1_275/A gnd OAI21X1_253/B vdd NAND2X1
XINVX1_500 INVX1_500/A gnd INVX1_500/Y vdd INVX1
XDFFPOSX1_318 AOI22X1_159/C CLKBUF1_51/Y OAI21X1_482/Y gnd vdd DFFPOSX1
XNOR2X1_135 gnd INVX1_369/Y gnd NOR2X1_135/Y vdd NOR2X1
XOAI21X1_102 AND2X2_2/Y NOR2X1_49/B INVX1_105/Y gnd OAI21X1_102/Y vdd OAI21X1
XXNOR2X1_45 BUFX2_117/Y BUFX2_77/Y gnd XNOR2X1_45/Y vdd XNOR2X1
XNAND2X1_216 INVX1_235/A INVX1_249/A gnd NAND2X1_216/Y vdd NAND2X1
XINVX1_464 INVX1_464/A gnd INVX1_464/Y vdd INVX1
XDFFPOSX1_282 AOI22X1_141/C CLKBUF1_17/Y OAI21X1_428/Y gnd vdd DFFPOSX1
XNAND2X1_180 NOR2X1_73/A BUFX2_67/Y gnd NAND2X1_181/B vdd NAND2X1
XDFFPOSX1_246 OAI21X1_373/C CLKBUF1_1/Y OAI21X1_374/Y gnd vdd DFFPOSX1
XAOI21X1_78 INVX1_541/Y AOI21X1_78/B AOI21X1_78/C gnd AOI21X1_78/Y vdd AOI21X1
XINVX1_428 BUFX2_116/Y gnd INVX1_428/Y vdd INVX1
XBUFX2_81 BUFX2_79/A gnd BUFX2_81/Y vdd BUFX2
XNAND2X1_144 BUFX2_72/Y INVX1_139/Y gnd OAI21X1_136/B vdd NAND2X1
XDFFPOSX1_210 OAI21X1_319/C CLKBUF1_36/Y OAI21X1_320/Y gnd vdd DFFPOSX1
XAOI21X1_42 INVX1_289/Y AOI21X1_42/B AOI21X1_42/C gnd AOI21X1_42/Y vdd AOI21X1
XINVX1_392 INVX1_392/A gnd INVX1_392/Y vdd INVX1
XNAND2X1_108 INVX1_93/A NAND2X1_108/B gnd AOI22X1_31/A vdd NAND2X1
XBUFX2_45 BUFX2_44/A gnd INVX1_55/A vdd BUFX2
XDFFPOSX1_174 AOI22X1_87/C CLKBUF1_22/Y OAI21X1_265/Y gnd vdd DFFPOSX1
XOAI21X1_90 INVX1_83/A INVX1_90/Y OAI21X1_89/Y gnd OAI21X1_90/Y vdd OAI21X1
XAOI22X1_176 INVX1_602/A INVX1_601/Y INVX1_603/Y AOI22X1_176/D gnd AOI22X1_176/Y vdd
+ AOI22X1
XOAI21X1_535 INVX1_601/Y INVX1_604/Y OAI21X1_535/C gnd OAI21X1_536/C vdd OAI21X1
XINVX1_356 BUFX2_122/Y gnd INVX1_356/Y vdd INVX1
XAOI22X1_83 AOI22X1_83/A AND2X2_68/Y AOI22X1_83/C NOR2X1_101/Y gnd AOI22X1_83/Y vdd
+ AOI22X1
XNAND2X1_69 INVX1_44/A NAND2X1_68/Y gnd AOI22X1_17/A vdd NAND2X1
XDFFPOSX1_72 INVX1_107/A CLKBUF1_15/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 AOI22X1_69/C CLKBUF1_45/Y OAI21X1_209/Y gnd vdd DFFPOSX1
XAOI22X1_140 INVX1_476/A INVX1_475/Y INVX1_477/Y AOI22X1_140/D gnd OAI21X1_430/B vdd
+ AOI22X1
XOAI21X1_54 INVX1_48/Y INVX1_51/Y AOI22X1_19/C gnd OAI21X1_55/C vdd OAI21X1
XOAI21X1_499 INVX1_559/Y INVX1_562/Y OAI21X1_499/C gnd OAI21X1_499/Y vdd OAI21X1
XINVX1_320 BUFX2_30/Y gnd INVX1_320/Y vdd INVX1
XAOI22X1_47 AOI22X1_47/A AND2X2_47/Y AOI22X1_47/C NOR2X1_62/Y gnd AOI22X1_47/Y vdd
+ AOI22X1
XOAI21X1_18 NOR2X1_18/Y AOI21X1_2/Y INVX1_6/A gnd OAI21X1_18/Y vdd OAI21X1
XDFFPOSX1_36 INVX1_44/A CLKBUF1_24/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XNAND2X1_33 request_put[4] NOR2X1_17/Y gnd NAND2X1_33/Y vdd NAND2X1
XINVX1_284 INVX1_284/A gnd INVX1_284/Y vdd INVX1
XAOI22X1_104 NAND2X1_7/A INVX1_349/Y INVX1_351/Y AOI22X1_104/D gnd AOI22X1_104/Y vdd
+ AOI22X1
XDFFPOSX1_102 AOI22X1_51/C CLKBUF1_30/Y OAI21X1_154/Y gnd vdd DFFPOSX1
XOAI21X1_463 INVX1_517/Y INVX1_520/Y AOI22X1_153/C gnd OAI21X1_463/Y vdd OAI21X1
XAOI22X1_11 INVX1_34/A AOI22X1_9/B OR2X2_4/A AOI22X1_9/D gnd AOI22X1_11/Y vdd AOI22X1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_427 INVX1_475/Y INVX1_478/Y AOI22X1_141/C gnd OAI21X1_427/Y vdd OAI21X1
XINVX1_248 AND2X2_63/B gnd INVX1_248/Y vdd INVX1
XNAND3X1_74 AND2X2_6/Y NOR2X1_88/B INVX1_233/Y gnd NAND3X1_74/Y vdd NAND3X1
XFILL_24_1 gnd vdd FILL
XINVX1_212 NAND2X1_9/B gnd INVX1_212/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XNAND3X1_38 AND2X2_2/Y NOR2X1_49/B INVX1_107/Y gnd NAND3X1_39/B vdd NAND3X1
XOAI21X1_391 INVX1_433/Y INVX1_436/Y AOI22X1_129/C gnd OAI21X1_392/C vdd OAI21X1
XFILL_14_2_1 gnd vdd FILL
XNAND2X1_505 INVX1_588/A BUFX2_12/Y gnd NAND2X1_506/B vdd NAND2X1
XFILL_16_0_0 gnd vdd FILL
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XAND2X2_107 INVX1_473/A INVX1_466/A gnd NOR2X1_178/B vdd AND2X2
XINVX1_176 INVX1_167/A gnd NOR2X1_71/B vdd INVX1
XOAI21X1_355 INVX1_391/Y INVX1_394/Y AOI22X1_117/C gnd OAI21X1_355/Y vdd OAI21X1
XNAND2X1_469 BUFX2_75/Y INVX1_548/A gnd NAND2X1_469/Y vdd NAND2X1
XFILL_2_0_2 gnd vdd FILL
XAND2X2_80 AND2X2_80/A AND2X2_79/B gnd AND2X2_80/Y vdd AND2X2
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XOAI21X1_319 INVX1_349/Y INVX1_352/Y OAI21X1_319/C gnd OAI21X1_319/Y vdd OAI21X1
XNAND2X1_433 INVX1_513/A INVX1_506/A gnd NOR3X1_6/A vdd NAND2X1
XAND2X2_44 INVX1_125/A INVX1_129/A gnd AND2X2_44/Y vdd AND2X2
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd BUFX2_65/A vdd NOR3X1
XINVX1_104 AND2X2_2/Y gnd INVX1_104/Y vdd INVX1
XOAI21X1_283 INVX1_311/Y NAND2X1_279/Y OAI21X1_283/C gnd OAI21X1_283/Y vdd OAI21X1
XNAND2X1_397 BUFX2_114/Y INVX1_457/Y gnd NAND2X1_397/Y vdd NAND2X1
XAOI22X1_2 INVX1_20/A AOI22X1_4/B request_put[1] AOI22X1_4/D gnd AOI22X1_2/Y vdd AOI22X1
XFILL_23_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_83 gnd INVX1_215/Y gnd NOR2X1_83/Y vdd NOR2X1
XFILL_21_2_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_247 INVX1_266/Y NAND2X1_246/Y NOR2X1_98/Y gnd AOI21X1_39/C vdd OAI21X1
XNAND2X1_361 AND2X2_5/A NAND2X1_361/B gnd NAND2X1_361/Y vdd NAND2X1
XFILL_11_3 gnd vdd FILL
XINVX1_609 INVX1_609/A gnd INVX1_609/Y vdd INVX1
XFILL_9_0_2 gnd vdd FILL
XNOR2X1_47 INVX1_98/A INVX1_99/Y gnd NOR2X1_47/Y vdd NOR2X1
XOAI21X1_211 INVX1_228/Y AOI22X1_68/Y AOI22X1_69/Y gnd OAI21X1_211/Y vdd OAI21X1
XNOR2X1_244 INVX1_623/A INVX1_624/Y gnd NOR2X1_244/Y vdd NOR2X1
XNAND2X1_325 AND2X2_2/Y INVX1_363/Y gnd OAI21X1_333/B vdd NAND2X1
XCLKBUF1_35 BUFX2_5/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XINVX1_573 BUFX2_124/Y gnd INVX1_573/Y vdd INVX1
XNAND3X1_157 NOR2X1_201/Y NAND3X1_156/Y OAI21X1_462/Y gnd NAND3X1_157/Y vdd NAND3X1
XOAI21X1_175 INVX1_193/A INVX1_207/A INVX1_200/A gnd NAND2X1_183/B vdd OAI21X1
XXNOR2X1_2 INVX1_43/A INVX1_41/A gnd AOI21X1_7/B vdd XNOR2X1
XNOR2X1_11 NOR2X1_11/A NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_208 INVX1_539/A INVX1_540/Y gnd NOR2X1_208/Y vdd NOR2X1
XNAND2X1_289 AND2X2_12/B BUFX2_19/Y gnd NAND2X1_289/Y vdd NAND2X1
XDFFPOSX1_355 INVX1_606/A CLKBUF1_32/Y OAI21X1_538/Y gnd vdd DFFPOSX1
XBUFX2_122 NOR3X1_2/Y gnd BUFX2_122/Y vdd BUFX2
XINVX1_537 BUFX2_32/Y gnd INVX1_537/Y vdd INVX1
XNAND3X1_121 NOR2X1_147/Y NAND3X1_121/B NAND3X1_121/C gnd NAND3X1_121/Y vdd NAND3X1
XOAI21X1_139 AND2X2_5/Y NOR2X1_62/B INVX1_147/Y gnd OAI21X1_139/Y vdd OAI21X1
XNOR2X1_172 INVX1_455/A INVX1_456/Y gnd NOR2X1_172/Y vdd NOR2X1
XXNOR2X1_82 BUFX2_11/Y INVX1_601/A gnd XNOR2X1_82/Y vdd XNOR2X1
XFILL_28_2_1 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XNAND2X1_253 BUFX2_58/Y INVX1_272/Y gnd OAI21X1_254/B vdd NAND2X1
XINVX1_501 INVX1_501/A gnd INVX1_501/Y vdd INVX1
XDFFPOSX1_319 INVX1_283/A CLKBUF1_22/Y OAI21X1_484/Y gnd vdd DFFPOSX1
XXNOR2X1_46 BUFX2_118/Y BUFX2_84/Y gnd AOI21X1_51/B vdd XNOR2X1
XNOR2X1_136 INVX1_371/A INVX1_372/Y gnd NOR2X1_136/Y vdd NOR2X1
XNAND2X1_217 NAND2X1_216/Y OAI21X1_212/Y gnd AND2X2_60/B vdd NAND2X1
XOAI21X1_103 INVX1_106/A INVX1_104/Y OAI21X1_102/Y gnd NAND3X1_39/C vdd OAI21X1
XDFFPOSX1_283 INVX1_480/A CLKBUF1_17/Y OAI21X1_430/Y gnd vdd DFFPOSX1
XINVX1_465 INVX1_430/A gnd INVX1_465/Y vdd INVX1
XXNOR2X1_10 INVX1_99/A INVX1_97/A gnd XNOR2X1_10/Y vdd XNOR2X1
XNAND2X1_181 INVX1_184/A NAND2X1_181/B gnd AOI22X1_57/A vdd NAND2X1
XNOR2X1_100 gnd INVX1_271/Y gnd NOR2X1_100/Y vdd NOR2X1
XINVX1_429 INVX1_429/A gnd INVX1_429/Y vdd INVX1
XDFFPOSX1_247 INVX1_417/A CLKBUF1_8/Y OAI21X1_376/Y gnd vdd DFFPOSX1
XAOI21X1_79 INVX1_548/Y AOI21X1_79/B AOI21X1_79/C gnd AOI21X1_79/Y vdd AOI21X1
XBUFX2_82 BUFX2_79/A gnd BUFX2_82/Y vdd BUFX2
XNAND2X1_145 BUFX2_46/Y INVX1_142/Y gnd AOI22X1_44/D vdd NAND2X1
XDFFPOSX1_211 INVX1_354/A CLKBUF1_36/Y OAI21X1_322/Y gnd vdd DFFPOSX1
XAOI21X1_43 INVX1_296/Y AOI21X1_43/B AOI21X1_43/C gnd AOI21X1_43/Y vdd AOI21X1
XINVX1_393 BUFX2_36/Y gnd INVX1_393/Y vdd INVX1
XBUFX2_46 BUFX2_47/A gnd BUFX2_46/Y vdd BUFX2
XNAND2X1_109 INVX1_97/A INVX1_100/A gnd OAI21X1_98/B vdd NAND2X1
XDFFPOSX1_175 INVX1_291/A CLKBUF1_22/Y OAI21X1_267/Y gnd vdd DFFPOSX1
XOAI21X1_91 INVX1_90/Y INVX1_93/Y AOI22X1_31/C gnd OAI21X1_92/C vdd OAI21X1
XAOI22X1_177 AOI22X1_177/A AND2X2_137/Y OAI21X1_535/C NOR2X1_238/Y gnd OAI21X1_538/C
+ vdd AOI22X1
XOAI21X1_536 INVX1_605/Y OAI21X1_536/B OAI21X1_536/C gnd OAI21X1_536/Y vdd OAI21X1
XINVX1_357 INVX1_357/A gnd INVX1_357/Y vdd INVX1
XAOI22X1_84 INVX1_280/A INVX1_279/Y INVX1_281/Y AOI22X1_84/D gnd AOI22X1_84/Y vdd
+ AOI22X1
XBUFX2_10 BUFX2_8/A gnd BUFX2_10/Y vdd BUFX2
XOAI21X1_55 INVX1_52/Y NAND2X1_70/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XNAND2X1_70 BUFX2_56/Y INVX1_51/A gnd NAND2X1_70/Y vdd NAND2X1
XDFFPOSX1_73 AND2X2_2/B CLKBUF1_43/Y NAND3X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 OR2X2_4/B CLKBUF1_45/Y OAI21X1_211/Y gnd vdd DFFPOSX1
XAOI22X1_141 NAND2X1_417/Y AND2X2_110/Y AOI22X1_141/C NOR2X1_184/Y gnd OAI21X1_430/C
+ vdd AOI22X1
XOAI21X1_500 INVX1_563/Y NAND2X1_479/Y OAI21X1_499/Y gnd OAI21X1_500/Y vdd OAI21X1
XINVX1_321 INVX1_582/A gnd INVX1_321/Y vdd INVX1
XAOI22X1_48 AND2X2_7/B INVX1_153/Y INVX1_155/Y AOI22X1_48/D gnd AOI22X1_48/Y vdd AOI22X1
XDFFPOSX1_103 INVX1_165/A CLKBUF1_27/Y OAI21X1_156/Y gnd vdd DFFPOSX1
XOAI21X1_19 INVX1_15/Y OR2X2_1/B OAI21X1_19/C gnd AOI22X1_4/D vdd OAI21X1
XDFFPOSX1_37 INVX1_42/A CLKBUF1_24/Y NAND3X1_21/Y gnd vdd DFFPOSX1
XNAND2X1_34 request_put[5] NOR2X1_17/Y gnd OAI21X1_15/C vdd NAND2X1
XAOI22X1_105 AOI22X1_105/A AND2X2_83/Y OAI21X1_319/C NOR2X1_130/Y gnd AOI22X1_105/Y
+ vdd AOI22X1
XOAI21X1_464 INVX1_521/Y NAND2X1_446/Y OAI21X1_463/Y gnd OAI21X1_464/Y vdd OAI21X1
XINVX1_285 BUFX2_32/Y gnd INVX1_285/Y vdd INVX1
XAOI22X1_12 INVX1_35/A AOI22X1_9/B OR2X2_4/B AOI22X1_9/D gnd NAND2X1_57/B vdd AOI22X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XNAND3X1_75 NOR2X1_87/Y NAND3X1_74/Y NAND3X1_75/C gnd NAND3X1_75/Y vdd NAND3X1
XOAI21X1_428 INVX1_479/Y NAND2X1_413/Y OAI21X1_427/Y gnd OAI21X1_428/Y vdd OAI21X1
XFILL_24_2 gnd vdd FILL
XOAI21X1_392 INVX1_437/Y NAND2X1_380/Y OAI21X1_392/C gnd OAI21X1_392/Y vdd OAI21X1
XINVX1_213 INVX1_221/A gnd INVX1_213/Y vdd INVX1
XINVX1_95 INVX1_87/A gnd INVX1_95/Y vdd INVX1
XFILL_16_0_1 gnd vdd FILL
XNAND3X1_39 NOR2X1_48/Y NAND3X1_39/B NAND3X1_39/C gnd NAND3X1_39/Y vdd NAND3X1
XFILL_14_2_2 gnd vdd FILL
XNAND2X1_506 INVX1_590/A NAND2X1_506/B gnd AOI22X1_173/A vdd NAND2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XAND2X2_108 BUFX2_84/Y INVX1_430/A gnd AND2X2_108/Y vdd AND2X2
XINVX1_177 AND2X2_50/B gnd INVX1_177/Y vdd INVX1
XOAI21X1_356 INVX1_395/Y NAND2X1_347/Y OAI21X1_355/Y gnd OAI21X1_356/Y vdd OAI21X1
XNAND2X1_470 INVX1_547/A INVX1_545/Y gnd NAND2X1_470/Y vdd NAND2X1
XAND2X2_81 BUFX2_22/Y INVX1_46/A gnd AND2X2_81/Y vdd AND2X2
XINVX1_141 BUFX2_72/Y gnd INVX1_141/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XOAI21X1_320 INVX1_353/Y OAI21X1_320/B OAI21X1_319/Y gnd OAI21X1_320/Y vdd OAI21X1
XNAND2X1_434 INVX1_525/A INVX1_520/A gnd NOR3X1_6/B vdd NAND2X1
XFILL_15_3_0 gnd vdd FILL
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XAND2X2_45 BUFX2_50/Y OAI21X1_3/Y gnd AND2X2_45/Y vdd AND2X2
XINVX1_105 AND2X2_2/B gnd INVX1_105/Y vdd INVX1
XOAI21X1_284 INVX1_308/Y NAND2X1_280/Y NOR2X1_111/Y gnd AOI21X1_45/C vdd OAI21X1
XNAND2X1_398 INVX1_455/A AND2X2_9/Y gnd NAND2X1_399/B vdd NAND2X1
XAOI22X1_3 INVX1_21/A AOI22X1_4/B request_put[2] AOI22X1_4/D gnd AOI22X1_3/Y vdd AOI22X1
XFILL_23_0_1 gnd vdd FILL
XFILL_1_3_2 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_84 INVX1_217/A INVX1_218/Y gnd NOR2X1_84/Y vdd NOR2X1
XFILL_21_2_2 gnd vdd FILL
XOAI21X1_248 INVX1_270/Y AOI22X1_80/Y AOI22X1_81/Y gnd OAI21X1_248/Y vdd OAI21X1
XNAND2X1_362 BUFX2_40/Y AND2X2_6/A gnd OAI21X1_374/B vdd NAND2X1
XINVX1_610 INVX1_76/A gnd INVX1_610/Y vdd INVX1
XNOR2X1_48 gnd INVX1_103/Y gnd NOR2X1_48/Y vdd NOR2X1
XOAI21X1_212 INVX1_235/A INVX1_249/A INVX1_242/A gnd OAI21X1_212/Y vdd OAI21X1
XNAND2X1_326 INVX1_363/A INVX1_366/Y gnd NAND2X1_326/Y vdd NAND2X1
XCLKBUF1_36 BUFX2_1/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XXNOR2X1_3 INVX1_41/A BUFX2_56/Y gnd XNOR2X1_3/Y vdd XNOR2X1
XNAND3X1_158 BUFX2_66/Y INVX1_526/Y INVX1_527/Y gnd NAND3X1_159/B vdd NAND3X1
XINVX1_574 INVX1_574/A gnd INVX1_574/Y vdd INVX1
XOAI21X1_176 AND2X2_3/Y NOR2X1_75/B INVX1_189/Y gnd OAI21X1_176/Y vdd OAI21X1
XFILL_22_3_0 gnd vdd FILL
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd BUFX2_67/A vdd NOR2X1
XNOR2X1_209 INVX1_564/A INVX1_557/A gnd NOR2X1_210/A vdd NOR2X1
XNAND2X1_290 INVX1_317/A NAND2X1_289/Y gnd AOI22X1_95/A vdd NAND2X1
XNAND3X1_122 BUFX2_41/Y INVX1_400/Y INVX1_401/Y gnd NAND3X1_123/B vdd NAND3X1
XDFFPOSX1_356 INVX1_604/A CLKBUF1_32/Y AOI21X1_87/Y gnd vdd DFFPOSX1
XINVX1_538 BUFX2_64/Y gnd INVX1_538/Y vdd INVX1
XBUFX2_123 NOR3X1_7/Y gnd INVX1_566/A vdd BUFX2
XOAI21X1_140 BUFX2_47/Y INVX1_146/Y OAI21X1_139/Y gnd NAND3X1_51/C vdd OAI21X1
XNOR2X1_173 INVX1_480/A INVX1_473/A gnd NOR2X1_174/A vdd NOR2X1
XFILL_28_2_2 gnd vdd FILL
XXNOR2X1_83 INVX1_76/A BUFX2_9/Y gnd AOI21X1_88/B vdd XNOR2X1
XFILL_8_3_2 gnd vdd FILL
XNAND2X1_254 AND2X2_9/Y INVX1_275/Y gnd AOI22X1_82/D vdd NAND2X1
XDFFPOSX1_320 AND2X2_15/A CLKBUF1_22/Y AOI21X1_78/Y gnd vdd DFFPOSX1
XINVX1_502 INVX1_89/A gnd INVX1_502/Y vdd INVX1
XOAI21X1_104 INVX1_104/Y INVX1_107/Y AOI22X1_35/C gnd OAI21X1_105/C vdd OAI21X1
XXNOR2X1_47 AND2X2_1/Y BUFX2_122/Y gnd AOI21X1_52/B vdd XNOR2X1
XNAND2X1_218 AND2X2_6/Y INVX1_233/A gnd OAI21X1_216/B vdd NAND2X1
XNOR2X1_137 AND2X2_88/A AND2X2_87/B gnd NOR2X1_138/A vdd NOR2X1
XDFFPOSX1_284 INVX1_478/A CLKBUF1_42/Y AOI21X1_69/Y gnd vdd DFFPOSX1
XINVX1_466 INVX1_466/A gnd INVX1_466/Y vdd INVX1
XXNOR2X1_11 INVX1_106/A AND2X2_2/Y gnd AOI21X1_16/B vdd XNOR2X1
XFILL_15_1 gnd vdd FILL
XNOR2X1_101 AND2X2_9/B INVX1_274/Y gnd NOR2X1_101/Y vdd NOR2X1
XNAND2X1_182 INVX1_193/A INVX1_207/A gnd NAND2X1_182/Y vdd NAND2X1
XINVX1_430 INVX1_430/A gnd INVX1_430/Y vdd INVX1
XDFFPOSX1_248 AND2X2_6/A CLKBUF1_15/Y AOI21X1_60/Y gnd vdd DFFPOSX1
XAOI21X1_80 INVX1_555/Y AOI21X1_80/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XBUFX2_83 BUFX2_85/A gnd BUFX2_83/Y vdd BUFX2
XNAND2X1_146 INVX1_140/A BUFX2_72/Y gnd NAND2X1_146/Y vdd NAND2X1
XDFFPOSX1_212 INVX1_352/A CLKBUF1_33/Y AOI21X1_51/Y gnd vdd DFFPOSX1
XAOI21X1_44 INVX1_303/Y XNOR2X1_39/Y AOI21X1_44/C gnd AOI21X1_44/Y vdd AOI21X1
XINVX1_394 INVX1_394/A gnd INVX1_394/Y vdd INVX1
XBUFX2_47 BUFX2_47/A gnd BUFX2_47/Y vdd BUFX2
XNAND2X1_110 INVX1_99/A INVX1_97/Y gnd OAI21X1_99/B vdd NAND2X1
XDFFPOSX1_176 INVX1_289/A CLKBUF1_22/Y AOI21X1_42/Y gnd vdd DFFPOSX1
XOAI21X1_92 INVX1_94/Y OAI21X1_92/B OAI21X1_92/C gnd OAI21X1_92/Y vdd OAI21X1
XAOI22X1_178 INVX1_609/A INVX1_608/Y INVX1_610/Y AOI22X1_178/D gnd AOI22X1_178/Y vdd
+ AOI22X1
XOAI21X1_537 INVX1_602/Y NAND2X1_513/Y NOR2X1_237/Y gnd AOI21X1_87/C vdd OAI21X1
XINVX1_358 AND2X2_1/Y gnd INVX1_358/Y vdd INVX1
XAOI22X1_85 AOI22X1_85/A AND2X2_69/Y AOI22X1_85/C AOI22X1_85/D gnd AOI22X1_85/Y vdd
+ AOI22X1
XBUFX2_11 BUFX2_8/A gnd BUFX2_11/Y vdd BUFX2
XDFFPOSX1_74 AOI22X1_37/C CLKBUF1_39/Y DFFPOSX1_74/D gnd vdd DFFPOSX1
XOAI21X1_56 INVX1_49/Y NAND2X1_71/Y NOR2X1_31/Y gnd AOI21X1_8/C vdd OAI21X1
XNAND2X1_71 INVX1_41/A INVX1_48/Y gnd NAND2X1_71/Y vdd NAND2X1
XAOI22X1_142 INVX1_483/A INVX1_482/Y INVX1_484/Y NAND2X1_420/Y gnd AOI22X1_142/Y vdd
+ AOI22X1
XDFFPOSX1_140 INVX1_226/A CLKBUF1_45/Y AOI21X1_33/Y gnd vdd DFFPOSX1
XOAI21X1_501 INVX1_560/Y OAI21X1_501/B NOR2X1_219/Y gnd AOI21X1_81/C vdd OAI21X1
XINVX1_322 AND2X2_18/B gnd INVX1_322/Y vdd INVX1
XAOI22X1_49 AOI22X1_49/A AND2X2_48/Y AOI22X1_49/C NOR2X1_64/Y gnd AOI22X1_49/Y vdd
+ AOI22X1
XNAND2X1_35 request_put[6] NOR2X1_17/Y gnd OAI21X1_16/C vdd NAND2X1
XDFFPOSX1_104 INVX1_163/A CLKBUF1_30/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XOAI21X1_20 NOR2X1_18/Y AOI21X1_2/Y INVX1_8/A gnd OAI21X1_20/Y vdd OAI21X1
XDFFPOSX1_38 AOI22X1_19/C CLKBUF1_12/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XINVX1_286 INVX1_575/A gnd INVX1_286/Y vdd INVX1
XAOI22X1_106 INVX1_357/A INVX1_356/Y INVX1_358/Y NAND2X1_321/Y gnd AOI22X1_106/Y vdd
+ AOI22X1
XOAI21X1_465 INVX1_518/Y OAI21X1_465/B NOR2X1_201/Y gnd AOI21X1_75/C vdd OAI21X1
XAOI22X1_13 INVX1_36/A AOI22X1_9/B INVX1_39/A AOI22X1_9/D gnd AOI22X1_13/Y vdd AOI22X1
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_429 INVX1_476/Y NAND2X1_414/Y NOR2X1_183/Y gnd AOI21X1_69/C vdd OAI21X1
XFILL_10_1_0 gnd vdd FILL
XINVX1_250 BUFX2_31/Y gnd INVX1_250/Y vdd INVX1
XNAND3X1_76 INVX1_237/A INVX1_239/Y INVX1_240/Y gnd NAND3X1_76/Y vdd NAND3X1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XOAI21X1_393 INVX1_434/Y NAND2X1_381/Y NOR2X1_165/Y gnd AOI21X1_63/C vdd OAI21X1
XINVX1_214 INVX1_395/A gnd INVX1_214/Y vdd INVX1
XFILL_16_0_2 gnd vdd FILL
XNAND3X1_40 AND2X2_4/Y NOR2X1_51/B INVX1_114/Y gnd NAND3X1_41/B vdd NAND3X1
XNAND2X1_507 BUFX2_78/Y INVX1_597/A gnd NAND2X1_507/Y vdd NAND2X1
XINVX1_60 OR2X2_5/A gnd INVX1_60/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XAND2X2_109 BUFX2_91/Y INVX1_395/A gnd AND2X2_109/Y vdd AND2X2
XOAI21X1_357 INVX1_392/Y OAI21X1_357/B NOR2X1_147/Y gnd AOI21X1_57/C vdd OAI21X1
XNAND2X1_471 BUFX2_74/Y INVX1_548/Y gnd AOI22X1_160/D vdd NAND2X1
XAND2X2_82 BUFX2_73/Y INVX1_88/A gnd AND2X2_82/Y vdd AND2X2
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XOAI21X1_321 INVX1_350/Y NAND2X1_315/Y NOR2X1_129/Y gnd AOI21X1_51/C vdd OAI21X1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XNAND2X1_435 INVX1_539/A INVX1_532/A gnd NOR3X1_6/C vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XAND2X2_46 BUFX2_46/Y AND2X2_46/B gnd AND2X2_46/Y vdd AND2X2
XFILL_15_3_1 gnd vdd FILL
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd BUFX2_8/A vdd NOR3X1
XINVX1_106 INVX1_106/A gnd NOR2X1_49/B vdd INVX1
XOAI21X1_285 INVX1_312/Y AOI22X1_92/Y AOI22X1_93/Y gnd OAI21X1_285/Y vdd OAI21X1
XNAND2X1_399 AND2X2_9/A NAND2X1_399/B gnd AOI22X1_135/A vdd NAND2X1
XAOI22X1_4 INVX1_22/A AOI22X1_4/B request_put[3] AOI22X1_4/D gnd AOI22X1_4/Y vdd AOI22X1
XAND2X2_10 INVX1_485/A AND2X2_10/B gnd INVX1_484/A vdd AND2X2
XFILL_23_0_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XNOR2X1_85 gnd INVX1_222/Y gnd NOR2X1_85/Y vdd NOR2X1
XNAND2X1_363 AND2X2_6/Y INVX1_412/Y gnd OAI21X1_375/B vdd NAND2X1
XOAI21X1_249 INVX1_277/A INVX1_291/A INVX1_284/A gnd NAND2X1_251/B vdd OAI21X1
XINVX1_611 INVX1_611/A gnd INVX1_611/Y vdd INVX1
XNOR2X1_49 AND2X2_2/B NOR2X1_49/B gnd NOR2X1_49/Y vdd NOR2X1
XOAI21X1_213 AND2X2_6/Y NOR2X1_88/B INVX1_231/Y gnd OAI21X1_213/Y vdd OAI21X1
XNAND2X1_327 INVX1_364/A AND2X2_2/Y gnd NAND2X1_328/B vdd NAND2X1
XNAND3X1_159 NOR2X1_203/Y NAND3X1_159/B OAI21X1_468/Y gnd NAND3X1_159/Y vdd NAND3X1
XCLKBUF1_37 BUFX2_6/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XFILL_24_1_0 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XXNOR2X1_4 BUFX2_69/Y INVX1_55/A gnd AOI21X1_9/B vdd XNOR2X1
XINVX1_575 INVX1_575/A gnd INVX1_575/Y vdd INVX1
XNOR2X1_13 INVX1_1/A NOR2X1_11/B gnd NOR2X1_13/Y vdd NOR2X1
XOAI21X1_177 INVX1_204/A INVX1_188/Y OAI21X1_176/Y gnd NAND3X1_63/C vdd OAI21X1
XFILL_4_2_0 gnd vdd FILL
XNOR2X1_210 NOR2X1_210/A NOR2X1_210/B gnd INVX1_570/A vdd NOR2X1
XNAND2X1_291 INVX1_582/A INVX1_324/A gnd NAND2X1_291/Y vdd NAND2X1
XNAND3X1_123 NOR2X1_149/Y NAND3X1_123/B NAND3X1_123/C gnd NAND3X1_123/Y vdd NAND3X1
XDFFPOSX1_357 INVX1_602/A CLKBUF1_23/Y NAND3X1_181/Y gnd vdd DFFPOSX1
XBUFX2_124 NOR3X1_7/Y gnd BUFX2_124/Y vdd BUFX2
XINVX1_539 INVX1_539/A gnd INVX1_539/Y vdd INVX1
XOAI21X1_141 INVX1_146/Y INVX1_149/Y AOI22X1_47/C gnd OAI21X1_141/Y vdd OAI21X1
XXNOR2X1_84 INVX1_160/A BUFX2_8/Y gnd XNOR2X1_84/Y vdd XNOR2X1
XNOR2X1_174 NOR2X1_174/A NOR2X1_174/B gnd INVX1_486/A vdd NOR2X1
XNAND2X1_255 AND2X2_9/B BUFX2_58/Y gnd NAND2X1_255/Y vdd NAND2X1
XDFFPOSX1_321 INVX1_539/A CLKBUF1_51/Y NAND3X1_163/Y gnd vdd DFFPOSX1
XINVX1_503 INVX1_43/A gnd INVX1_503/Y vdd INVX1
XOAI21X1_105 INVX1_108/Y OAI21X1_105/B OAI21X1_105/C gnd DFFPOSX1_70/D vdd OAI21X1
XXNOR2X1_48 AND2X2_2/Y INVX1_363/A gnd AOI21X1_53/B vdd XNOR2X1
XNAND2X1_219 BUFX2_14/Y INVX1_230/Y gnd NAND2X1_219/Y vdd NAND2X1
XNOR2X1_138 NOR2X1_138/A AND2X2_87/Y gnd INVX1_402/A vdd NOR2X1
XDFFPOSX1_285 INVX1_476/A CLKBUF1_17/Y NAND3X1_145/Y gnd vdd DFFPOSX1
XINVX1_467 BUFX2_32/Y gnd INVX1_467/Y vdd INVX1
XXNOR2X1_12 INVX1_113/A AND2X2_4/Y gnd AOI21X1_17/B vdd XNOR2X1
XFILL_15_2 gnd vdd FILL
XNOR2X1_102 gnd INVX1_278/Y gnd NAND3X1_89/A vdd NOR2X1
XNAND2X1_183 NAND2X1_182/Y NAND2X1_183/B gnd AND2X2_53/B vdd NAND2X1
XINVX1_431 INVX1_431/A gnd INVX1_431/Y vdd INVX1
XDFFPOSX1_249 INVX1_413/A CLKBUF1_8/Y NAND3X1_127/Y gnd vdd DFFPOSX1
XAOI21X1_81 INVX1_562/Y AOI21X1_81/B AOI21X1_81/C gnd AOI21X1_81/Y vdd AOI21X1
XBUFX2_84 BUFX2_85/A gnd BUFX2_84/Y vdd BUFX2
XNAND2X1_147 INVX1_142/A NAND2X1_146/Y gnd AOI22X1_45/A vdd NAND2X1
XDFFPOSX1_213 NAND2X1_7/A CLKBUF1_33/Y NAND3X1_109/Y gnd vdd DFFPOSX1
XAOI21X1_45 INVX1_310/Y AOI21X1_45/B AOI21X1_45/C gnd AOI21X1_45/Y vdd AOI21X1
XINVX1_395 INVX1_395/A gnd INVX1_395/Y vdd INVX1
XBUFX2_48 BUFX2_47/A gnd BUFX2_48/Y vdd BUFX2
XNAND2X1_111 INVX1_97/A INVX1_100/Y gnd AOI22X1_32/D vdd NAND2X1
XOAI21X1_93 INVX1_91/Y OAI21X1_93/B NOR2X1_44/Y gnd AOI21X1_14/C vdd OAI21X1
XOAI21X1_538 INVX1_606/Y AOI22X1_176/Y OAI21X1_538/C gnd OAI21X1_538/Y vdd OAI21X1
XDFFPOSX1_177 AND2X2_17/B CLKBUF1_22/Y NAND3X1_91/Y gnd vdd DFFPOSX1
XAOI22X1_179 NAND2X1_521/Y AND2X2_138/Y AOI22X1_179/C NOR2X1_240/Y gnd AOI22X1_179/Y
+ vdd AOI22X1
XINVX1_359 AND2X2_1/A gnd INVX1_359/Y vdd INVX1
XBUFX2_12 BUFX2_8/A gnd BUFX2_12/Y vdd BUFX2
XAOI22X1_86 AND2X2_17/B INVX1_286/Y INVX1_288/Y AOI22X1_86/D gnd AOI22X1_86/Y vdd
+ AOI22X1
XDFFPOSX1_141 INVX1_224/A CLKBUF1_35/Y NAND3X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 INVX1_116/A CLKBUF1_1/Y OAI21X1_113/Y gnd vdd DFFPOSX1
XOAI21X1_57 INVX1_53/Y OAI21X1_57/B AOI22X1_19/Y gnd OAI21X1_57/Y vdd OAI21X1
XNAND2X1_72 BUFX2_56/Y INVX1_51/Y gnd NAND2X1_72/Y vdd NAND2X1
XAOI22X1_143 NAND2X1_422/Y AND2X2_111/Y OAI21X1_433/C NOR2X1_186/Y gnd AOI22X1_143/Y
+ vdd AOI22X1
XOAI21X1_502 INVX1_564/Y OAI21X1_502/B OAI21X1_502/C gnd OAI21X1_502/Y vdd OAI21X1
XINVX1_323 BUFX2_19/Y gnd INVX1_323/Y vdd INVX1
XAOI22X1_50 INVX1_161/A INVX1_160/Y INVX1_162/Y AOI22X1_50/D gnd AOI22X1_50/Y vdd
+ AOI22X1
XNAND2X1_36 INVX1_3/Y INVX1_15/Y gnd AND2X2_23/B vdd NAND2X1
XDFFPOSX1_105 INVX1_161/A CLKBUF1_30/Y NAND3X1_55/Y gnd vdd DFFPOSX1
XAOI22X1_107 AOI22X1_107/A AND2X2_84/Y OAI21X1_325/C NOR2X1_132/Y gnd AOI22X1_107/Y
+ vdd AOI22X1
XOAI21X1_21 NOR2X1_18/Y AOI21X1_2/Y INVX1_9/A gnd OAI21X1_21/Y vdd OAI21X1
XDFFPOSX1_39 INVX1_45/A CLKBUF1_24/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XINVX1_287 AND2X2_17/B gnd INVX1_287/Y vdd INVX1
XOAI21X1_466 INVX1_522/Y AOI22X1_152/Y AOI22X1_153/Y gnd OAI21X1_466/Y vdd OAI21X1
XAOI22X1_14 INVX1_37/A AOI22X1_9/B INVX1_38/A AOI22X1_9/D gnd AOI22X1_14/Y vdd AOI22X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XOAI21X1_430 INVX1_480/Y OAI21X1_430/B OAI21X1_430/C gnd OAI21X1_430/Y vdd OAI21X1
XFILL_10_1_1 gnd vdd FILL
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XNAND3X1_77 NOR2X1_89/Y NAND3X1_76/Y NAND3X1_77/C gnd NAND3X1_77/Y vdd NAND3X1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XOAI21X1_394 INVX1_438/Y OAI21X1_394/B OAI21X1_394/C gnd OAI21X1_394/Y vdd OAI21X1
XINVX1_215 INVX1_89/A gnd INVX1_215/Y vdd INVX1
XNAND3X1_41 NOR2X1_50/Y NAND3X1_41/B NAND3X1_41/C gnd NAND3X1_41/Y vdd NAND3X1
XNAND2X1_508 BUFX2_13/Y INVX1_594/Y gnd NAND2X1_508/Y vdd NAND2X1
XINVX1_179 INVX1_171/A gnd INVX1_179/Y vdd INVX1
XINVX1_61 BUFX2_32/Y gnd INVX1_61/Y vdd INVX1
XAND2X2_110 INVX1_475/A INVX1_479/A gnd AND2X2_110/Y vdd AND2X2
XNAND2X1_472 NAND2X1_4/A INVX1_547/A gnd NAND2X1_472/Y vdd NAND2X1
XOAI21X1_358 INVX1_396/Y OAI21X1_358/B OAI21X1_358/C gnd OAI21X1_358/Y vdd OAI21X1
XAND2X2_83 BUFX2_86/Y INVX1_430/A gnd AND2X2_83/Y vdd AND2X2
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_143 AND2X2_46/B gnd INVX1_143/Y vdd INVX1
XOAI21X1_322 INVX1_354/Y AOI22X1_104/Y AOI22X1_105/Y gnd OAI21X1_322/Y vdd OAI21X1
XNAND2X1_436 BUFX2_25/Y INVX1_506/A gnd NAND2X1_436/Y vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAND2X2_47 AND2X2_5/Y AND2X2_47/B gnd AND2X2_47/Y vdd AND2X2
XFILL_15_3_2 gnd vdd FILL
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XOAI21X1_286 INVX1_319/A INVX1_333/A INVX1_326/A gnd OAI21X1_286/Y vdd OAI21X1
XNAND2X1_400 INVX1_471/A INVX1_464/A gnd NOR3X1_5/A vdd NAND2X1
XAOI22X1_5 INVX1_23/A AOI22X1_4/B request_put[4] AOI22X1_4/D gnd AOI22X1_5/Y vdd AOI22X1
XAND2X2_11 AND2X2_11/A NOR2X1_90/A gnd INVX1_237/A vdd AND2X2
XNOR2X1_86 INVX1_224/A INVX1_225/Y gnd NOR2X1_86/Y vdd NOR2X1
XOAI21X1_250 AND2X2_9/Y INVX1_274/Y INVX1_273/Y gnd OAI21X1_251/C vdd OAI21X1
XNAND2X1_364 BUFX2_40/Y INVX1_415/Y gnd NAND2X1_364/Y vdd NAND2X1
XFILL_28_1 gnd vdd FILL
XNOR2X1_50 gnd INVX1_110/Y gnd NOR2X1_50/Y vdd NOR2X1
XINVX1_612 INVX1_612/A gnd INVX1_612/Y vdd INVX1
XOAI21X1_214 BUFX2_14/Y INVX1_230/Y OAI21X1_213/Y gnd NAND3X1_75/C vdd OAI21X1
XNAND2X1_328 AND2X2_2/A NAND2X1_328/B gnd AOI22X1_109/A vdd NAND2X1
XNAND3X1_160 BUFX2_62/Y INVX1_533/Y INVX1_534/Y gnd NAND3X1_161/B vdd NAND3X1
XINVX1_576 INVX1_576/A gnd INVX1_576/Y vdd INVX1
XCLKBUF1_38 BUFX2_6/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XFILL_6_0_0 gnd vdd FILL
XFILL_24_1_1 gnd vdd FILL
XXNOR2X1_5 INVX1_64/A AND2X2_1/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_22_3_2 gnd vdd FILL
XNOR2X1_14 NOR2X1_9/B NOR2X1_11/A gnd NOR2X1_14/Y vdd NOR2X1
XOAI21X1_178 INVX1_188/Y INVX1_191/Y AOI22X1_59/C gnd OAI21X1_179/C vdd OAI21X1
XFILL_4_2_1 gnd vdd FILL
XNOR2X1_211 INVX1_564/A INVX1_550/A gnd NOR2X1_211/Y vdd NOR2X1
XNAND2X1_292 BUFX2_19/Y INVX1_321/Y gnd NAND2X1_292/Y vdd NAND2X1
XNAND3X1_124 BUFX2_39/Y INVX1_407/Y INVX1_408/Y gnd NAND3X1_124/Y vdd NAND3X1
XBUFX2_125 NOR3X1_7/Y gnd BUFX2_125/Y vdd BUFX2
XINVX1_540 INVX1_279/A gnd INVX1_540/Y vdd INVX1
XDFFPOSX1_358 AOI22X1_179/C CLKBUF1_9/Y OAI21X1_542/Y gnd vdd DFFPOSX1
XOAI21X1_142 INVX1_150/Y NAND2X1_150/Y OAI21X1_141/Y gnd OAI21X1_142/Y vdd OAI21X1
XXNOR2X1_85 INVX1_624/A BUFX2_12/Y gnd XNOR2X1_85/Y vdd XNOR2X1
XNOR2X1_175 INVX1_480/A INVX1_466/A gnd NOR2X1_176/A vdd NOR2X1
XNAND2X1_256 INVX1_275/A NAND2X1_255/Y gnd AOI22X1_83/A vdd NAND2X1
XDFFPOSX1_322 AOI22X1_161/C CLKBUF1_48/Y OAI21X1_488/Y gnd vdd DFFPOSX1
XINVX1_504 NAND2X1_2/B gnd INVX1_504/Y vdd INVX1
XXNOR2X1_49 AND2X2_3/Y INVX1_370/A gnd XNOR2X1_49/Y vdd XNOR2X1
XOAI21X1_106 INVX1_105/Y OAI21X1_106/B NOR2X1_48/Y gnd AOI21X1_16/C vdd OAI21X1
XNOR2X1_139 AND2X2_88/A AND2X2_88/B gnd NOR2X1_140/A vdd NOR2X1
XNAND2X1_220 AND2X2_6/Y INVX1_233/Y gnd AOI22X1_70/D vdd NAND2X1
XDFFPOSX1_286 OAI21X1_433/C CLKBUF1_4/Y OAI21X1_434/Y gnd vdd DFFPOSX1
XINVX1_468 BUFX2_91/Y gnd INVX1_468/Y vdd INVX1
XXNOR2X1_13 INVX1_113/A AND2X2_42/A gnd AOI21X1_18/B vdd XNOR2X1
XFILL_15_3 gnd vdd FILL
XNAND2X1_184 AND2X2_3/Y INVX1_191/A gnd OAI21X1_179/B vdd NAND2X1
XNOR2X1_103 INVX1_280/A INVX1_281/Y gnd AOI22X1_85/D vdd NOR2X1
XDFFPOSX1_250 OAI21X1_379/C CLKBUF1_8/Y OAI21X1_380/Y gnd vdd DFFPOSX1
XAOI21X1_82 INVX1_569/Y XNOR2X1_77/Y AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XINVX1_432 BUFX2_31/Y gnd INVX1_432/Y vdd INVX1
XBUFX2_85 BUFX2_85/A gnd BUFX2_85/Y vdd BUFX2
XNAND2X1_148 INVX1_151/A INVX1_165/A gnd NAND2X1_148/Y vdd NAND2X1
XDFFPOSX1_214 OAI21X1_325/C CLKBUF1_32/Y OAI21X1_326/Y gnd vdd DFFPOSX1
XINVX1_396 AND2X2_88/A gnd INVX1_396/Y vdd INVX1
XAOI21X1_46 INVX1_317/Y XNOR2X1_41/Y AOI21X1_46/C gnd AOI21X1_46/Y vdd AOI21X1
XBUFX2_49 BUFX2_47/A gnd BUFX2_49/Y vdd BUFX2
XNAND2X1_112 INVX1_98/A BUFX2_72/Y gnd NAND2X1_112/Y vdd NAND2X1
XOAI21X1_94 INVX1_95/Y OAI21X1_94/B OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XAOI22X1_180 INVX1_616/A INVX1_615/Y INVX1_617/Y AOI22X1_180/D gnd OAI21X1_550/B vdd
+ AOI22X1
XDFFPOSX1_178 AOI22X1_89/C CLKBUF1_37/Y OAI21X1_271/Y gnd vdd DFFPOSX1
XINVX1_360 AND2X2_84/B gnd INVX1_360/Y vdd INVX1
XAOI21X1_10 INVX1_65/Y XNOR2X1_5/Y AOI21X1_10/C gnd AOI21X1_10/Y vdd AOI21X1
XOAI21X1_539 BUFX2_9/Y INVX1_610/Y INVX1_609/Y gnd OAI21X1_539/Y vdd OAI21X1
XBUFX2_13 BUFX2_8/A gnd BUFX2_13/Y vdd BUFX2
XNAND2X1_73 INVX1_4/A INVX1_41/A gnd NAND2X1_74/B vdd NAND2X1
XAOI22X1_87 AOI22X1_87/A AND2X2_70/Y AOI22X1_87/C NOR2X1_105/Y gnd AOI22X1_87/Y vdd
+ AOI22X1
XDFFPOSX1_142 AOI22X1_71/C CLKBUF1_31/Y OAI21X1_216/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 INVX1_114/A CLKBUF1_39/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XOAI21X1_58 INVX1_55/A INVX1_57/Y INVX1_56/Y gnd OAI21X1_59/C vdd OAI21X1
XAOI22X1_144 INVX1_490/A INVX1_489/Y INVX1_491/Y AOI22X1_144/D gnd OAI21X1_442/B vdd
+ AOI22X1
XOAI21X1_503 INVX1_566/A INVX1_568/Y INVX1_567/Y gnd OAI21X1_504/C vdd OAI21X1
XINVX1_324 INVX1_324/A gnd INVX1_324/Y vdd INVX1
XAOI22X1_51 AOI22X1_51/A AND2X2_49/Y AOI22X1_51/C NOR2X1_66/Y gnd AOI22X1_51/Y vdd
+ AOI22X1
XOAI21X1_22 NOR2X1_18/Y AOI21X1_2/Y INVX1_10/A gnd NAND2X1_40/A vdd OAI21X1
XNAND2X1_37 OAI21X1_18/Y AOI22X1_1/Y gnd NAND2X1_37/Y vdd NAND2X1
XDFFPOSX1_106 AOI22X1_53/C CLKBUF1_4/Y OAI21X1_160/Y gnd vdd DFFPOSX1
XAOI22X1_108 INVX1_364/A INVX1_363/Y INVX1_365/Y NAND2X1_326/Y gnd AOI22X1_108/Y vdd
+ AOI22X1
XINVX1_288 BUFX2_57/Y gnd INVX1_288/Y vdd INVX1
XDFFPOSX1_40 INVX1_51/A CLKBUF1_24/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XOAI21X1_467 BUFX2_66/Y INVX1_526/Y INVX1_525/Y gnd OAI21X1_468/C vdd OAI21X1
XAOI22X1_15 NOR2X1_27/Y INVX1_38/Y OAI21X1_45/Y NAND3X1_19/Y gnd NAND3X1_17/A vdd
+ AOI22X1
XFILL_10_1_2 gnd vdd FILL
XOAI21X1_431 BUFX2_134/Y INVX1_484/Y INVX1_483/Y gnd OAI21X1_431/Y vdd OAI21X1
XINVX1_252 NOR2X1_95/A gnd INVX1_252/Y vdd INVX1
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XNAND3X1_78 INVX1_244/A NOR2X1_92/B INVX1_247/Y gnd NAND3X1_79/B vdd NAND3X1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XOAI21X1_395 INVX1_440/A INVX1_442/Y INVX1_441/Y gnd OAI21X1_395/Y vdd OAI21X1
XNAND3X1_42 AND2X2_42/A NOR2X1_53/B INVX1_121/Y gnd NAND3X1_42/Y vdd NAND3X1
XINVX1_216 BUFX2_55/Y gnd INVX1_216/Y vdd INVX1
XNAND2X1_509 BUFX2_78/Y INVX1_597/Y gnd NAND2X1_509/Y vdd NAND2X1
XAND2X2_111 BUFX2_129/Y INVX1_486/A gnd AND2X2_111/Y vdd AND2X2
XINVX1_180 BUFX2_31/Y gnd NOR2X1_72/B vdd INVX1
XOAI21X1_359 BUFX2_41/Y INVX1_400/Y INVX1_399/Y gnd OAI21X1_360/C vdd OAI21X1
XCLKBUF1_1 BUFX2_3/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XINVX1_62 AND2X2_1/Y gnd INVX1_62/Y vdd INVX1
XFILL_11_2_0 gnd vdd FILL
XNAND2X1_473 INVX1_548/A NAND2X1_472/Y gnd AOI22X1_161/A vdd NAND2X1
XAND2X2_84 AND2X2_85/A AND2X2_84/B gnd AND2X2_84/Y vdd AND2X2
XINVX1_26 BUFX2_31/Y gnd INVX1_26/Y vdd INVX1
XINVX1_144 OR2X2_3/B gnd INVX1_144/Y vdd INVX1
XOAI21X1_323 BUFX2_122/Y INVX1_358/Y INVX1_357/Y gnd OAI21X1_323/Y vdd OAI21X1
XNAND2X1_437 BUFX2_61/Y INVX1_503/Y gnd NAND2X1_437/Y vdd NAND2X1
XFILL_17_1_2 gnd vdd FILL
XAND2X2_48 AND2X2_7/Y INVX1_157/A gnd AND2X2_48/Y vdd AND2X2
XINVX1_108 INVX1_368/A gnd INVX1_108/Y vdd INVX1
XNAND2X1_401 INVX1_483/A INVX1_478/A gnd NOR3X1_5/B vdd NAND2X1
XAOI22X1_6 INVX1_24/A AOI22X1_4/B request_put[5] AOI22X1_4/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_287 INVX1_498/A INVX1_316/Y INVX1_315/Y gnd OAI21X1_287/Y vdd OAI21X1
XFILL_6_1 gnd vdd FILL
XAND2X2_12 INVX1_499/A AND2X2_12/B gnd INVX1_498/A vdd AND2X2
XNOR2X1_87 gnd NOR2X1_87/B gnd NOR2X1_87/Y vdd NOR2X1
XOAI21X1_251 BUFX2_58/Y INVX1_272/Y OAI21X1_251/C gnd NAND3X1_87/C vdd OAI21X1
XNAND2X1_365 INVX1_413/A AND2X2_6/Y gnd NAND2X1_366/B vdd NAND2X1
XFILL_28_2 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XNOR2X1_51 AND2X2_4/B NOR2X1_51/B gnd NOR2X1_51/Y vdd NOR2X1
XINVX1_613 INVX1_80/A gnd INVX1_613/Y vdd INVX1
XOAI21X1_215 INVX1_230/Y INVX1_233/Y AOI22X1_71/C gnd OAI21X1_216/C vdd OAI21X1
XNAND2X1_329 INVX1_370/A AND2X2_3/A gnd NAND2X1_329/Y vdd NAND2X1
XCLKBUF1_39 BUFX2_3/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XFILL_24_1_2 gnd vdd FILL
XNAND3X1_161 NOR2X1_205/Y NAND3X1_161/B OAI21X1_474/Y gnd NAND3X1_161/Y vdd NAND3X1
XINVX1_577 INVX1_577/A gnd INVX1_577/Y vdd INVX1
XOAI21X1_179 INVX1_192/Y OAI21X1_179/B OAI21X1_179/C gnd OAI21X1_179/Y vdd OAI21X1
XFILL_4_2_2 gnd vdd FILL
XFILL_6_0_1 gnd vdd FILL
XXNOR2X1_6 BUFX2_43/Y INVX1_69/A gnd XNOR2X1_6/Y vdd XNOR2X1
XNOR2X1_15 NOR3X1_1/B NOR3X1_1/C gnd NAND3X1_8/C vdd NOR2X1
XNOR2X1_212 NOR2X1_211/Y AND2X2_124/Y gnd INVX1_577/A vdd NOR2X1
XNAND2X1_293 INVX1_582/A INVX1_324/Y gnd AOI22X1_96/D vdd NAND2X1
XDFFPOSX1_359 INVX1_80/A CLKBUF1_9/Y OAI21X1_544/Y gnd vdd DFFPOSX1
XNAND3X1_125 NOR2X1_151/Y NAND3X1_124/Y OAI21X1_366/Y gnd NAND3X1_125/Y vdd NAND3X1
XBUFX2_126 NOR3X1_7/Y gnd INVX1_554/A vdd BUFX2
XINVX1_541 AND2X2_15/A gnd INVX1_541/Y vdd INVX1
XOAI21X1_143 INVX1_147/Y NAND2X1_151/Y NOR2X1_61/Y gnd AOI21X1_22/C vdd OAI21X1
XNOR2X1_176 NOR2X1_176/A NOR2X1_176/B gnd INVX1_493/A vdd NOR2X1
XNAND2X1_257 INVX1_279/A INVX1_282/A gnd NAND2X1_257/Y vdd NAND2X1
XDFFPOSX1_323 INVX1_550/A CLKBUF1_19/Y OAI21X1_490/Y gnd vdd DFFPOSX1
XINVX1_505 BUFX2_61/Y gnd INVX1_505/Y vdd INVX1
XOAI21X1_107 INVX1_109/Y AOI22X1_34/Y AOI22X1_35/Y gnd OAI21X1_107/Y vdd OAI21X1
XNOR2X1_140 NOR2X1_140/A AND2X2_88/Y gnd INVX1_409/A vdd NOR2X1
XXNOR2X1_50 BUFX2_36/Y BUFX2_75/Y gnd AOI21X1_55/B vdd XNOR2X1
XFILL_25_2_0 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XNAND2X1_221 AND2X2_6/B BUFX2_14/Y gnd NAND2X1_222/B vdd NAND2X1
XDFFPOSX1_287 INVX1_487/A CLKBUF1_31/Y OAI21X1_436/Y gnd vdd DFFPOSX1
XINVX1_469 INVX1_469/A gnd INVX1_469/Y vdd INVX1
XXNOR2X1_14 BUFX2_82/Y INVX1_125/A gnd AOI21X1_19/B vdd XNOR2X1
XNAND2X1_185 INVX1_190/A INVX1_188/Y gnd NAND2X1_185/Y vdd NAND2X1
XNOR2X1_104 gnd INVX1_285/Y gnd NOR2X1_104/Y vdd NOR2X1
XDFFPOSX1_251 AND2X2_98/B CLKBUF1_36/Y OAI21X1_382/Y gnd vdd DFFPOSX1
XAOI21X1_83 INVX1_576/Y XNOR2X1_78/Y AOI21X1_83/C gnd AOI21X1_83/Y vdd AOI21X1
XINVX1_433 BUFX2_96/Y gnd INVX1_433/Y vdd INVX1
XBUFX2_86 BUFX2_85/A gnd BUFX2_86/Y vdd BUFX2
XNAND2X1_149 NAND2X1_148/Y OAI21X1_138/Y gnd AND2X2_46/B vdd NAND2X1
XINVX1_397 BUFX2_35/Y gnd INVX1_397/Y vdd INVX1
XAOI21X1_47 INVX1_324/Y XNOR2X1_42/Y AOI21X1_47/C gnd AOI21X1_47/Y vdd AOI21X1
XDFFPOSX1_215 INVX1_66/A CLKBUF1_9/Y OAI21X1_328/Y gnd vdd DFFPOSX1
XBUFX2_50 BUFX2_54/A gnd BUFX2_50/Y vdd BUFX2
XNAND2X1_113 INVX1_100/A NAND2X1_112/Y gnd AOI22X1_33/A vdd NAND2X1
XOAI21X1_95 INVX1_97/A INVX1_99/Y INVX1_98/Y gnd OAI21X1_95/Y vdd OAI21X1
XDFFPOSX1_179 INVX1_479/A CLKBUF1_37/Y OAI21X1_273/Y gnd vdd DFFPOSX1
XAOI22X1_181 NAND2X1_526/Y AND2X2_139/Y AOI22X1_181/C NOR2X1_242/Y gnd OAI21X1_550/C
+ vdd AOI22X1
XAOI21X1_11 INVX1_72/Y XNOR2X1_6/Y OAI21X1_75/Y gnd AOI21X1_11/Y vdd AOI21X1
XOAI21X1_540 INVX1_76/A INVX1_608/Y OAI21X1_539/Y gnd NAND3X1_183/C vdd OAI21X1
XINVX1_361 INVX1_66/A gnd INVX1_361/Y vdd INVX1
XBUFX2_14 BUFX2_17/A gnd BUFX2_14/Y vdd BUFX2
XAOI22X1_88 INVX1_294/A INVX1_293/Y INVX1_295/Y AOI22X1_88/D gnd AOI22X1_88/Y vdd
+ AOI22X1
XNAND2X1_74 INVX1_51/A NAND2X1_74/B gnd AOI22X1_19/A vdd NAND2X1
XAOI22X1_145 AOI22X1_145/A AND2X2_112/Y AOI22X1_145/C NOR2X1_188/Y gnd AOI22X1_145/Y
+ vdd AOI22X1
XDFFPOSX1_143 INVX1_235/A CLKBUF1_31/Y OAI21X1_218/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 AND2X2_4/B CLKBUF1_15/Y NAND3X1_41/Y gnd vdd DFFPOSX1
XOAI21X1_59 BUFX2_68/Y INVX1_55/Y OAI21X1_59/C gnd NAND3X1_25/C vdd OAI21X1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XOAI21X1_504 AND2X2_42/A INVX1_566/Y OAI21X1_504/C gnd NAND3X1_171/C vdd OAI21X1
XAOI22X1_52 INVX1_168/A INVX1_167/Y INVX1_169/Y AOI22X1_52/D gnd AOI22X1_52/Y vdd
+ AOI22X1
XOAI21X1_23 NOR2X1_18/Y AOI21X1_2/Y INVX1_11/A gnd OAI21X1_23/Y vdd OAI21X1
XNAND2X1_38 OAI21X1_20/Y AOI22X1_2/Y gnd NAND2X1_38/Y vdd NAND2X1
XDFFPOSX1_41 INVX1_4/A CLKBUF1_12/Y NAND3X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 INVX1_430/A CLKBUF1_33/Y OAI21X1_162/Y gnd vdd DFFPOSX1
XAOI22X1_109 AOI22X1_109/A AND2X2_85/Y OAI21X1_331/C NOR2X1_134/Y gnd OAI21X1_334/C
+ vdd AOI22X1
XOAI21X1_468 INVX1_69/A INVX1_524/Y OAI21X1_468/C gnd OAI21X1_468/Y vdd OAI21X1
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XFILL_19_1 gnd vdd FILL
XAOI22X1_16 INVX1_42/A INVX1_41/Y INVX1_43/Y AOI22X1_16/D gnd OAI21X1_51/B vdd AOI22X1
XOAI21X1_432 INVX1_484/A INVX1_482/Y OAI21X1_431/Y gnd OAI21X1_432/Y vdd OAI21X1
XINVX1_253 BUFX2_95/Y gnd INVX1_253/Y vdd INVX1
XNAND3X1_79 NOR2X1_91/Y NAND3X1_79/B NAND3X1_79/C gnd NAND3X1_79/Y vdd NAND3X1
XOAI21X1_396 AND2X2_7/Y INVX1_440/Y OAI21X1_395/Y gnd OAI21X1_396/Y vdd OAI21X1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XNAND3X1_43 NOR2X1_52/Y NAND3X1_42/Y NAND3X1_43/C gnd NAND3X1_43/Y vdd NAND3X1
XNAND2X1_510 NAND2X1_6/B BUFX2_13/Y gnd NAND2X1_511/B vdd NAND2X1
XINVX1_63 AND2X2_1/B gnd INVX1_63/Y vdd INVX1
XINVX1_181 BUFX2_108/Y gnd INVX1_181/Y vdd INVX1
XAND2X2_112 BUFX2_129/Y INVX1_493/A gnd AND2X2_112/Y vdd AND2X2
XOAI21X1_360 AND2X2_4/Y INVX1_398/Y OAI21X1_360/C gnd NAND3X1_123/C vdd OAI21X1
XFILL_11_2_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XCLKBUF1_2 BUFX2_7/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XNAND2X1_474 BUFX2_94/Y INVX1_555/A gnd OAI21X1_494/B vdd NAND2X1
XAND2X2_85 AND2X2_85/A INVX1_367/A gnd AND2X2_85/Y vdd AND2X2
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_145 BUFX2_35/Y gnd NOR2X1_61/B vdd INVX1
XOAI21X1_324 AND2X2_1/Y INVX1_356/Y OAI21X1_323/Y gnd OAI21X1_324/Y vdd OAI21X1
XNAND2X1_438 BUFX2_25/Y INVX1_506/Y gnd AOI22X1_148/D vdd NAND2X1
XAND2X2_49 INVX1_160/A AND2X2_49/B gnd AND2X2_49/Y vdd AND2X2
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XOAI21X1_288 BUFX2_18/Y INVX1_314/Y OAI21X1_287/Y gnd NAND3X1_99/C vdd OAI21X1
XNAND2X1_402 INVX1_497/A INVX1_490/A gnd NOR3X1_5/C vdd NAND2X1
XAOI22X1_7 INVX1_25/A AOI22X1_4/B request_put[6] AOI22X1_4/D gnd AOI22X1_7/Y vdd AOI22X1
XAND2X2_13 AND2X2_13/A INVX1_70/A gnd INVX1_69/A vdd AND2X2
XNOR2X1_88 AND2X2_6/B NOR2X1_88/B gnd NOR2X1_88/Y vdd NOR2X1
XOAI21X1_252 INVX1_272/Y INVX1_275/Y AOI22X1_83/C gnd OAI21X1_253/C vdd OAI21X1
XNAND2X1_366 AND2X2_6/A NAND2X1_366/B gnd AOI22X1_123/A vdd NAND2X1
XFILL_20_0_0 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XINVX1_614 BUFX2_35/Y gnd INVX1_614/Y vdd INVX1
XFILL_18_2_1 gnd vdd FILL
XNOR2X1_52 gnd NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XNAND2X1_330 AND2X2_3/Y INVX1_370/Y gnd OAI21X1_339/B vdd NAND2X1
XOAI21X1_216 INVX1_234/Y OAI21X1_216/B OAI21X1_216/C gnd OAI21X1_216/Y vdd OAI21X1
XNAND3X1_162 BUFX2_64/Y INVX1_540/Y INVX1_541/Y gnd NAND3X1_162/Y vdd NAND3X1
XINVX1_578 INVX1_578/A gnd INVX1_578/Y vdd INVX1
XCLKBUF1_40 BUFX2_2/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XOAI21X1_180 INVX1_189/Y NAND2X1_185/Y NOR2X1_74/Y gnd AOI21X1_28/C vdd OAI21X1
XFILL_6_0_2 gnd vdd FILL
XNOR2X1_16 gnd INVX1_14/Y gnd NOR2X1_16/Y vdd NOR2X1
XXNOR2X1_7 BUFX2_42/Y INVX1_76/A gnd XNOR2X1_7/Y vdd XNOR2X1
XNOR2X1_213 INVX1_557/A INVX1_550/A gnd NOR2X1_213/Y vdd NOR2X1
XNAND2X1_294 AND2X2_18/B BUFX2_19/Y gnd NAND2X1_295/B vdd NAND2X1
XNAND3X1_126 BUFX2_40/Y INVX1_414/Y INVX1_415/Y gnd NAND3X1_126/Y vdd NAND3X1
XDFFPOSX1_360 INVX1_611/A CLKBUF1_9/Y AOI21X1_88/Y gnd vdd DFFPOSX1
XBUFX2_127 NOR3X1_7/Y gnd INVX1_547/A vdd BUFX2
XINVX1_542 INVX1_542/A gnd INVX1_542/Y vdd INVX1
XOAI21X1_144 INVX1_151/Y AOI22X1_46/Y AOI22X1_47/Y gnd OAI21X1_144/Y vdd OAI21X1
XNOR2X1_177 INVX1_473/A INVX1_466/A gnd NOR2X1_177/Y vdd NOR2X1
XNAND2X1_258 BUFX2_59/Y INVX1_279/Y gnd OAI21X1_260/B vdd NAND2X1
XDFFPOSX1_324 INVX1_548/A CLKBUF1_19/Y AOI21X1_79/Y gnd vdd DFFPOSX1
XINVX1_506 INVX1_506/A gnd INVX1_506/Y vdd INVX1
XOAI21X1_108 AND2X2_4/Y NOR2X1_51/B INVX1_112/Y gnd OAI21X1_108/Y vdd OAI21X1
XXNOR2X1_51 BUFX2_37/Y BUFX2_81/Y gnd AOI21X1_56/B vdd XNOR2X1
XFILL_27_0_0 gnd vdd FILL
XFILL_25_2_1 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XNAND2X1_222 INVX1_233/A NAND2X1_222/B gnd AOI22X1_71/A vdd NAND2X1
XFILL_7_1_0 gnd vdd FILL
XNOR2X1_141 AND2X2_87/B AND2X2_88/B gnd NOR2X1_141/Y vdd NOR2X1
XDFFPOSX1_288 INVX1_485/A CLKBUF1_4/Y AOI21X1_70/Y gnd vdd DFFPOSX1
XINVX1_470 BUFX2_132/Y gnd INVX1_470/Y vdd INVX1
XXNOR2X1_15 INVX1_125/A BUFX2_50/Y gnd AOI21X1_20/B vdd XNOR2X1
XNAND2X1_186 AND2X2_3/Y INVX1_191/Y gnd AOI22X1_58/D vdd NAND2X1
XNOR2X1_105 AND2X2_17/B INVX1_288/Y gnd NOR2X1_105/Y vdd NOR2X1
XDFFPOSX1_252 INVX1_422/A CLKBUF1_8/Y AOI21X1_61/Y gnd vdd DFFPOSX1
XINVX1_434 INVX1_434/A gnd INVX1_434/Y vdd INVX1
XAOI21X1_84 INVX1_583/Y XNOR2X1_79/Y AOI21X1_84/C gnd AOI21X1_84/Y vdd AOI21X1
XBUFX2_87 BUFX2_85/A gnd BUFX2_87/Y vdd BUFX2
XNAND2X1_150 AND2X2_5/Y INVX1_149/A gnd NAND2X1_150/Y vdd NAND2X1
XINVX1_398 BUFX2_41/Y gnd INVX1_398/Y vdd INVX1
XAOI21X1_48 INVX1_331/Y XNOR2X1_43/Y AOI21X1_48/C gnd AOI21X1_48/Y vdd AOI21X1
XDFFPOSX1_216 AND2X2_1/A CLKBUF1_32/Y AOI21X1_52/Y gnd vdd DFFPOSX1
XBUFX2_51 BUFX2_54/A gnd BUFX2_51/Y vdd BUFX2
XNAND2X1_114 INVX1_109/A INVX1_123/A gnd NAND2X1_114/Y vdd NAND2X1
XOAI21X1_1 INVX1_6/Y NOR3X1_1/Y NAND3X1_5/Y gnd INVX1_52/A vdd OAI21X1
XOAI21X1_96 INVX1_99/A INVX1_97/Y OAI21X1_95/Y gnd OAI21X1_96/Y vdd OAI21X1
XDFFPOSX1_180 INVX1_296/A CLKBUF1_13/Y AOI21X1_43/Y gnd vdd DFFPOSX1
XAOI21X1_12 INVX1_79/Y XNOR2X1_7/Y OAI21X1_81/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI22X1_182 INVX1_623/A INVX1_622/Y INVX1_624/Y AOI22X1_182/D gnd OAI21X1_556/B vdd
+ AOI22X1
XINVX1_362 BUFX2_35/Y gnd INVX1_362/Y vdd INVX1
XOAI21X1_541 INVX1_608/Y INVX1_611/Y AOI22X1_179/C gnd OAI21X1_542/C vdd OAI21X1
XBUFX2_15 BUFX2_17/A gnd BUFX2_15/Y vdd BUFX2
XAOI22X1_89 AOI22X1_89/A AND2X2_72/Y AOI22X1_89/C AOI22X1_89/D gnd AOI22X1_89/Y vdd
+ AOI22X1
XDFFPOSX1_78 AOI22X1_39/C CLKBUF1_8/Y DFFPOSX1_78/D gnd vdd DFFPOSX1
XNAND2X1_75 BUFX2_43/Y INVX1_58/A gnd NAND2X1_75/Y vdd NAND2X1
XOAI21X1_60 INVX1_55/Y INVX1_58/Y AOI22X1_21/C gnd OAI21X1_61/C vdd OAI21X1
XDFFPOSX1_144 INVX1_233/A CLKBUF1_31/Y AOI21X1_34/Y gnd vdd DFFPOSX1
XOAI21X1_505 INVX1_566/Y INVX1_569/Y AOI22X1_167/C gnd OAI21X1_505/Y vdd OAI21X1
XAOI22X1_146 INVX1_497/A INVX1_496/Y INVX1_498/Y AOI22X1_146/D gnd AOI22X1_146/Y vdd
+ AOI22X1
XINVX1_326 INVX1_326/A gnd INVX1_326/Y vdd INVX1
XAOI22X1_53 AOI22X1_53/A AND2X2_51/Y AOI22X1_53/C NOR2X1_69/Y gnd AOI22X1_53/Y vdd
+ AOI22X1
XDFFPOSX1_108 INVX1_170/A CLKBUF1_4/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XNAND2X1_39 OAI21X1_21/Y AOI22X1_3/Y gnd NAND2X1_39/Y vdd NAND2X1
XOAI21X1_24 NOR2X1_18/Y AOI21X1_2/Y INVX1_12/A gnd NAND2X1_42/A vdd OAI21X1
XDFFPOSX1_42 AOI22X1_21/C CLKBUF1_11/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XAOI22X1_110 INVX1_371/A INVX1_370/Y INVX1_372/Y NAND2X1_331/Y gnd AOI22X1_110/Y vdd
+ AOI22X1
XOAI21X1_469 INVX1_524/Y INVX1_527/Y AOI22X1_155/C gnd OAI21X1_470/C vdd OAI21X1
XINVX1_290 INVX1_578/A gnd INVX1_290/Y vdd INVX1
XFILL_19_2 gnd vdd FILL
XAOI22X1_17 AOI22X1_17/A AND2X2_30/Y AOI22X1_17/C NOR2X1_30/Y gnd OAI21X1_51/C vdd
+ AOI22X1
XOAI21X1_433 INVX1_482/Y INVX1_485/Y OAI21X1_433/C gnd OAI21X1_434/C vdd OAI21X1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XNAND3X1_80 INVX1_251/A INVX1_253/Y INVX1_254/Y gnd NAND3X1_81/B vdd NAND3X1
XOAI21X1_397 INVX1_440/Y INVX1_443/Y OAI21X1_397/C gnd OAI21X1_397/Y vdd OAI21X1
XINVX1_218 INVX1_209/A gnd INVX1_218/Y vdd INVX1
XNAND2X1_511 INVX1_597/A NAND2X1_511/B gnd NAND2X1_511/Y vdd NAND2X1
XNAND3X1_44 INVX1_125/A NOR2X1_56/B INVX1_128/Y gnd NAND3X1_44/Y vdd NAND3X1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_182 NOR2X1_73/A gnd INVX1_182/Y vdd INVX1
XOAI21X1_361 INVX1_398/Y INVX1_401/Y OAI21X1_361/C gnd OAI21X1_361/Y vdd OAI21X1
XFILL_11_2_2 gnd vdd FILL
XAND2X2_113 BUFX2_132/Y INVX1_500/A gnd AND2X2_113/Y vdd AND2X2
XFILL_13_0_1 gnd vdd FILL
XCLKBUF1_3 BUFX2_7/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XNAND2X1_475 BUFX2_125/Y INVX1_552/Y gnd NAND2X1_475/Y vdd NAND2X1
XAND2X2_86 INVX1_370/A AND2X2_86/B gnd AND2X2_86/Y vdd AND2X2
XINVX1_146 AND2X2_5/Y gnd INVX1_146/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XOAI21X1_325 INVX1_356/Y INVX1_359/Y OAI21X1_325/C gnd OAI21X1_326/C vdd OAI21X1
XNAND2X1_439 NAND2X1_2/B BUFX2_61/Y gnd NAND2X1_439/Y vdd NAND2X1
XAND2X2_50 INVX1_168/A AND2X2_50/B gnd INVX1_167/A vdd AND2X2
XINVX1_110 BUFX2_35/Y gnd INVX1_110/Y vdd INVX1
XOAI21X1_289 INVX1_314/Y INVX1_317/Y AOI22X1_95/C gnd OAI21X1_290/C vdd OAI21X1
XNAND2X1_403 BUFX2_83/Y INVX1_464/A gnd OAI21X1_416/B vdd NAND2X1
XFILL_12_3_0 gnd vdd FILL
XAOI22X1_8 INVX1_30/A AOI22X1_9/B OR2X2_5/A AOI22X1_9/D gnd AOI22X1_8/Y vdd AOI22X1
XAND2X2_14 AND2X2_14/A INVX1_245/A gnd INVX1_244/A vdd AND2X2
XNOR2X1_89 gnd INVX1_236/Y gnd NOR2X1_89/Y vdd NOR2X1
XOAI21X1_253 INVX1_276/Y OAI21X1_253/B OAI21X1_253/C gnd OAI21X1_253/Y vdd OAI21X1
XNAND2X1_367 INVX1_429/A INVX1_422/A gnd NOR3X1_4/A vdd NAND2X1
XFILL_20_0_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XINVX1_615 BUFX2_8/Y gnd INVX1_615/Y vdd INVX1
XFILL_18_2_2 gnd vdd FILL
XOAI21X1_217 INVX1_231/Y NAND2X1_219/Y NOR2X1_87/Y gnd AOI21X1_34/C vdd OAI21X1
XNOR2X1_53 NOR2X1_53/A NOR2X1_53/B gnd NOR2X1_53/Y vdd NOR2X1
XNAND2X1_331 INVX1_370/A INVX1_373/Y gnd NAND2X1_331/Y vdd NAND2X1
XCLKBUF1_41 BUFX2_3/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XINVX1_579 BUFX2_33/Y gnd INVX1_579/Y vdd INVX1
XNOR2X1_17 INVX1_15/Y INVX1_19/Y gnd NOR2X1_17/Y vdd NOR2X1
XNAND3X1_163 NOR2X1_207/Y NAND3X1_162/Y NAND3X1_163/C gnd NAND3X1_163/Y vdd NAND3X1
XXNOR2X1_8 BUFX2_76/Y INVX1_83/A gnd XNOR2X1_8/Y vdd XNOR2X1
XOAI21X1_181 INVX1_193/Y AOI22X1_58/Y AOI22X1_59/Y gnd OAI21X1_181/Y vdd OAI21X1
XNOR2X1_214 NOR2X1_213/Y AND2X2_125/Y gnd INVX1_584/A vdd NOR2X1
XNAND2X1_295 INVX1_324/A NAND2X1_295/B gnd AOI22X1_97/A vdd NAND2X1
XNAND3X1_127 NOR2X1_153/Y NAND3X1_126/Y OAI21X1_372/Y gnd NAND3X1_127/Y vdd NAND3X1
XBUFX2_128 NOR3X1_7/Y gnd INVX1_580/A vdd BUFX2
XINVX1_543 INVX1_283/A gnd INVX1_543/Y vdd INVX1
XDFFPOSX1_361 INVX1_609/A CLKBUF1_40/Y NAND3X1_183/Y gnd vdd DFFPOSX1
XFILL_19_3_0 gnd vdd FILL
XOAI21X1_145 AND2X2_7/Y INVX1_155/Y INVX1_154/Y gnd OAI21X1_145/Y vdd OAI21X1
XNOR2X1_178 NOR2X1_177/Y NOR2X1_178/B gnd INVX1_500/A vdd NOR2X1
XNAND2X1_259 INVX1_279/A INVX1_282/Y gnd AOI22X1_84/D vdd NAND2X1
XFILL_10_1 gnd vdd FILL
XDFFPOSX1_325 NAND2X1_4/A CLKBUF1_48/Y NAND3X1_165/Y gnd vdd DFFPOSX1
XINVX1_507 INVX1_46/A gnd INVX1_507/Y vdd INVX1
XOAI21X1_109 INVX1_113/A INVX1_111/Y OAI21X1_108/Y gnd NAND3X1_41/C vdd OAI21X1
XFILL_27_0_1 gnd vdd FILL
XFILL_25_2_2 gnd vdd FILL
XXNOR2X1_52 BUFX2_36/Y BUFX2_88/Y gnd AOI21X1_57/B vdd XNOR2X1
XNAND2X1_223 INVX1_237/A INVX1_240/A gnd OAI21X1_222/B vdd NAND2X1
XFILL_5_3_2 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XNOR2X1_142 NOR2X1_141/Y AND2X2_89/Y gnd INVX1_416/A vdd NOR2X1
XDFFPOSX1_289 INVX1_483/A CLKBUF1_4/Y NAND3X1_147/Y gnd vdd DFFPOSX1
XINVX1_471 INVX1_471/A gnd INVX1_471/Y vdd INVX1
XXNOR2X1_16 BUFX2_72/Y BUFX2_49/Y gnd XNOR2X1_16/Y vdd XNOR2X1
XNOR2X1_106 NOR2X1_106/A NOR2X1_106/B gnd BUFX2_18/A vdd NOR2X1
XNAND2X1_187 AND2X2_3/B INVX1_190/A gnd NAND2X1_188/B vdd NAND2X1
XDFFPOSX1_253 INVX1_420/A CLKBUF1_23/Y NAND3X1_129/Y gnd vdd DFFPOSX1
XINVX1_435 BUFX2_112/Y gnd INVX1_435/Y vdd INVX1
XAOI21X1_85 INVX1_590/Y AOI21X1_85/B AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XBUFX2_88 BUFX2_88/A gnd BUFX2_88/Y vdd BUFX2
XNAND2X1_151 BUFX2_47/Y INVX1_146/Y gnd NAND2X1_151/Y vdd NAND2X1
XFILL_26_3_0 gnd vdd FILL
XDFFPOSX1_217 INVX1_357/A CLKBUF1_9/Y NAND3X1_111/Y gnd vdd DFFPOSX1
XINVX1_399 INVX1_399/A gnd INVX1_399/Y vdd INVX1
XAOI21X1_49 INVX1_338/Y AOI21X1_49/B AOI21X1_49/C gnd AOI21X1_49/Y vdd AOI21X1
XBUFX2_52 BUFX2_54/A gnd BUFX2_52/Y vdd BUFX2
XNAND2X1_115 NAND2X1_114/Y OAI21X1_101/Y gnd AND2X2_39/B vdd NAND2X1
XOAI21X1_97 INVX1_97/Y INVX1_100/Y AOI22X1_33/C gnd OAI21X1_98/C vdd OAI21X1
XOAI21X1_2 INVX1_8/Y NOR3X1_1/Y NAND3X1_6/Y gnd INVX1_94/A vdd OAI21X1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XDFFPOSX1_181 INVX1_294/A CLKBUF1_20/Y NAND3X1_93/Y gnd vdd DFFPOSX1
XAOI22X1_183 NAND2X1_531/Y AND2X2_140/Y AOI22X1_183/C NOR2X1_244/Y gnd AOI22X1_183/Y
+ vdd AOI22X1
XAOI21X1_13 INVX1_86/Y XNOR2X1_8/Y OAI21X1_87/Y gnd AOI21X1_13/Y vdd AOI21X1
XOAI21X1_542 INVX1_612/Y NAND2X1_517/Y OAI21X1_542/C gnd OAI21X1_542/Y vdd OAI21X1
XBUFX2_16 BUFX2_17/A gnd BUFX2_16/Y vdd BUFX2
XAOI22X1_90 INVX1_301/A INVX1_300/Y INVX1_302/Y AOI22X1_90/D gnd AOI22X1_90/Y vdd
+ AOI22X1
XDFFPOSX1_79 INVX1_123/A CLKBUF1_1/Y DFFPOSX1_79/D gnd vdd DFFPOSX1
XOAI21X1_61 INVX1_59/Y NAND2X1_75/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XNAND2X1_76 BUFX2_69/Y INVX1_55/Y gnd NAND2X1_76/Y vdd NAND2X1
XDFFPOSX1_145 AND2X2_6/B CLKBUF1_17/Y NAND3X1_75/Y gnd vdd DFFPOSX1
XOAI21X1_506 INVX1_570/Y NAND2X1_484/Y OAI21X1_505/Y gnd OAI21X1_506/Y vdd OAI21X1
XAOI22X1_147 AOI22X1_147/A AND2X2_113/Y OAI21X1_445/C NOR2X1_190/Y gnd OAI21X1_448/C
+ vdd AOI22X1
XINVX1_327 INVX1_89/A gnd INVX1_327/Y vdd INVX1
XAOI22X1_54 NOR2X1_71/A INVX1_174/Y NOR2X1_71/B AOI22X1_54/D gnd AOI22X1_54/Y vdd
+ AOI22X1
XNAND2X1_40 NAND2X1_40/A AOI22X1_4/Y gnd NAND2X1_40/Y vdd NAND2X1
XDFFPOSX1_109 INVX1_168/A CLKBUF1_4/Y NAND3X1_57/Y gnd vdd DFFPOSX1
XOAI21X1_25 NOR2X1_18/Y AOI21X1_2/Y INVX1_13/A gnd NAND2X1_43/A vdd OAI21X1
XDFFPOSX1_43 OR2X2_5/A CLKBUF1_11/Y OAI21X1_63/Y gnd vdd DFFPOSX1
XAOI22X1_111 NAND2X1_333/Y AND2X2_86/Y OAI21X1_337/C NOR2X1_136/Y gnd OAI21X1_340/C
+ vdd AOI22X1
XOAI21X1_470 INVX1_528/Y NAND2X1_451/Y OAI21X1_470/C gnd OAI21X1_470/Y vdd OAI21X1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XFILL_19_3 gnd vdd FILL
XAOI22X1_18 INVX1_4/A INVX1_48/Y INVX1_50/Y NAND2X1_72/Y gnd OAI21X1_57/B vdd AOI22X1
XOAI21X1_434 INVX1_486/Y NAND2X1_418/Y OAI21X1_434/C gnd OAI21X1_434/Y vdd OAI21X1
XINVX1_255 AND2X2_65/B gnd INVX1_255/Y vdd INVX1
XNAND3X1_81 NOR2X1_94/Y NAND3X1_81/B NAND3X1_81/C gnd NAND3X1_81/Y vdd NAND3X1
XOAI21X1_398 INVX1_444/Y NAND2X1_385/Y OAI21X1_397/Y gnd OAI21X1_398/Y vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XNAND2X1_512 INVX1_601/A INVX1_604/A gnd OAI21X1_536/B vdd NAND2X1
XNAND3X1_45 NOR2X1_55/Y NAND3X1_44/Y NAND3X1_45/C gnd NAND3X1_45/Y vdd NAND3X1
XFILL_13_0_2 gnd vdd FILL
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XCLKBUF1_4 BUFX2_5/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XINVX1_183 BUFX2_67/Y gnd NOR2X1_73/B vdd INVX1
XOAI21X1_362 INVX1_402/Y OAI21X1_362/B OAI21X1_361/Y gnd OAI21X1_362/Y vdd OAI21X1
XAND2X2_114 INVX1_522/A INVX1_515/A gnd AND2X2_114/Y vdd AND2X2
XNAND2X1_476 BUFX2_97/Y INVX1_555/Y gnd NAND2X1_476/Y vdd NAND2X1
XAND2X2_87 AND2X2_88/A AND2X2_87/B gnd AND2X2_87/Y vdd AND2X2
XINVX1_147 AND2X2_5/B gnd INVX1_147/Y vdd INVX1
XINVX1_29 EN_response_get gnd INVX1_29/Y vdd INVX1
XOAI21X1_326 INVX1_360/Y OAI21X1_326/B OAI21X1_326/C gnd OAI21X1_326/Y vdd OAI21X1
XNAND2X1_440 INVX1_506/A NAND2X1_439/Y gnd AOI22X1_149/A vdd NAND2X1
XAND2X2_51 INVX1_167/A INVX1_171/A gnd AND2X2_51/Y vdd AND2X2
XINVX1_111 AND2X2_4/Y gnd INVX1_111/Y vdd INVX1
XOAI21X1_290 INVX1_318/Y OAI21X1_290/B OAI21X1_290/C gnd OAI21X1_290/Y vdd OAI21X1
XNAND2X1_404 INVX1_463/A INVX1_461/Y gnd OAI21X1_417/B vdd NAND2X1
XAOI22X1_9 INVX1_32/A AOI22X1_9/B AOI22X1_9/C AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XFILL_12_3_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XAND2X2_15 AND2X2_15/A INVX1_280/A gnd INVX1_279/A vdd AND2X2
XNOR2X1_90 NOR2X1_90/A INVX1_239/Y gnd NOR2X1_90/Y vdd NOR2X1
XNAND2X1_368 INVX1_441/A INVX1_436/A gnd NOR3X1_4/B vdd NAND2X1
XOAI21X1_254 INVX1_273/Y OAI21X1_254/B NOR2X1_100/Y gnd AOI21X1_40/C vdd OAI21X1
XFILL_20_0_2 gnd vdd FILL
XFILL_0_1_2 gnd vdd FILL
XINVX1_616 INVX1_616/A gnd INVX1_616/Y vdd INVX1
XNOR2X1_54 NOR2X1_54/A NOR2X1_54/B gnd BUFX2_47/A vdd NOR2X1
XOAI21X1_218 INVX1_235/Y AOI22X1_70/Y AOI22X1_71/Y gnd OAI21X1_218/Y vdd OAI21X1
XNAND2X1_332 INVX1_371/A AND2X2_3/Y gnd NAND2X1_332/Y vdd NAND2X1
XNAND3X1_164 BUFX2_74/Y INVX1_547/Y INVX1_548/Y gnd NAND3X1_164/Y vdd NAND3X1
XCLKBUF1_42 BUFX2_2/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XINVX1_580 INVX1_580/A gnd INVX1_580/Y vdd INVX1
XNOR2X1_18 EN_request_put INVX1_16/Y gnd NOR2X1_18/Y vdd NOR2X1
XXNOR2X1_9 INVX1_83/A BUFX2_53/Y gnd XNOR2X1_9/Y vdd XNOR2X1
XOAI21X1_182 AND2X2_8/Y NOR2X1_77/B INVX1_196/Y gnd OAI21X1_182/Y vdd OAI21X1
XNOR2X1_215 gnd INVX1_544/Y gnd NOR2X1_215/Y vdd NOR2X1
XNAND2X1_296 INVX1_624/A INVX1_331/A gnd NAND2X1_296/Y vdd NAND2X1
XBUFX2_129 NOR3X1_5/Y gnd BUFX2_129/Y vdd BUFX2
XNAND3X1_128 BUFX2_80/Y INVX1_421/Y INVX1_422/Y gnd NAND3X1_128/Y vdd NAND3X1
XDFFPOSX1_362 AOI22X1_181/C CLKBUF1_39/Y OAI21X1_548/Y gnd vdd DFFPOSX1
XINVX1_544 INVX1_96/A gnd INVX1_544/Y vdd INVX1
XFILL_21_1_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_146 BUFX2_49/Y INVX1_153/Y OAI21X1_145/Y gnd NAND3X1_53/C vdd OAI21X1
XFILL_19_3_1 gnd vdd FILL
XNOR2X1_179 gnd INVX1_460/Y gnd NOR2X1_179/Y vdd NOR2X1
XNAND2X1_260 INVX1_280/A BUFX2_59/Y gnd NAND2X1_261/B vdd NAND2X1
XFILL_10_2 gnd vdd FILL
XDFFPOSX1_326 OAI21X1_493/C CLKBUF1_17/Y OAI21X1_494/Y gnd vdd DFFPOSX1
XINVX1_508 INVX1_508/A gnd INVX1_508/Y vdd INVX1
XFILL_27_0_2 gnd vdd FILL
XFILL_7_1_2 gnd vdd FILL
XOAI21X1_110 INVX1_111/Y INVX1_114/Y AOI22X1_37/C gnd OAI21X1_111/C vdd OAI21X1
XXNOR2X1_53 AND2X2_4/Y BUFX2_41/Y gnd AOI21X1_58/B vdd XNOR2X1
XNAND2X1_224 BUFX2_17/Y INVX1_237/Y gnd OAI21X1_223/B vdd NAND2X1
XNOR2X1_143 gnd INVX1_376/Y gnd NOR2X1_143/Y vdd NOR2X1
XDFFPOSX1_290 AOI22X1_145/C CLKBUF1_42/Y OAI21X1_440/Y gnd vdd DFFPOSX1
XINVX1_472 INVX1_395/A gnd INVX1_472/Y vdd INVX1
XXNOR2X1_17 BUFX2_47/Y AND2X2_5/Y gnd XNOR2X1_17/Y vdd XNOR2X1
XNOR2X1_107 gnd INVX1_292/Y gnd NAND3X1_93/A vdd NOR2X1
XNAND2X1_188 INVX1_191/A NAND2X1_188/B gnd AOI22X1_59/A vdd NAND2X1
XDFFPOSX1_254 OAI21X1_385/C CLKBUF1_33/Y OAI21X1_386/Y gnd vdd DFFPOSX1
XINVX1_436 INVX1_436/A gnd INVX1_436/Y vdd INVX1
XAOI21X1_86 INVX1_597/Y XNOR2X1_81/Y AOI21X1_86/C gnd AOI21X1_86/Y vdd AOI21X1
XBUFX2_89 BUFX2_88/A gnd BUFX2_89/Y vdd BUFX2
XNAND2X1_152 AND2X2_5/Y INVX1_149/Y gnd AOI22X1_46/D vdd NAND2X1
XFILL_26_3_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XDFFPOSX1_218 OAI21X1_331/C CLKBUF1_27/Y OAI21X1_332/Y gnd vdd DFFPOSX1
XFILL_8_2_0 gnd vdd FILL
XAOI21X1_50 INVX1_345/Y XNOR2X1_45/Y AOI21X1_50/C gnd AOI21X1_50/Y vdd AOI21X1
XINVX1_400 AND2X2_4/Y gnd INVX1_400/Y vdd INVX1
XBUFX2_53 BUFX2_54/A gnd BUFX2_53/Y vdd BUFX2
XNAND2X1_116 AND2X2_2/Y INVX1_107/A gnd OAI21X1_105/B vdd NAND2X1
XOAI21X1_98 INVX1_101/Y OAI21X1_98/B OAI21X1_98/C gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_3 INVX1_9/Y NOR3X1_1/Y NAND3X1_7/Y gnd OAI21X1_3/Y vdd OAI21X1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XAOI21X1_14 INVX1_93/Y XNOR2X1_9/Y AOI21X1_14/C gnd AOI21X1_14/Y vdd AOI21X1
XOAI21X1_543 INVX1_609/Y OAI21X1_543/B NOR2X1_239/Y gnd AOI21X1_88/C vdd OAI21X1
XDFFPOSX1_182 AOI22X1_91/C CLKBUF1_11/Y OAI21X1_277/Y gnd vdd DFFPOSX1
XBUFX2_17 BUFX2_17/A gnd BUFX2_17/Y vdd BUFX2
XAOI22X1_91 AOI22X1_91/A AND2X2_73/Y AOI22X1_91/C AOI22X1_91/D gnd AOI22X1_91/Y vdd
+ AOI22X1
XDFFPOSX1_146 AOI22X1_73/C CLKBUF1_4/Y OAI21X1_222/Y gnd vdd DFFPOSX1
XDFFPOSX1_80 INVX1_121/A CLKBUF1_1/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XNAND2X1_77 INVX1_55/A INVX1_58/Y gnd AOI22X1_20/D vdd NAND2X1
XOAI21X1_62 INVX1_56/Y NAND2X1_76/Y NOR2X1_33/Y gnd AOI21X1_9/C vdd OAI21X1
XOAI21X1_507 INVX1_567/Y OAI21X1_507/B NOR2X1_221/Y gnd AOI21X1_82/C vdd OAI21X1
XAOI22X1_148 NAND2X1_2/B INVX1_503/Y INVX1_505/Y AOI22X1_148/D gnd AOI22X1_148/Y vdd
+ AOI22X1
XINVX1_328 INVX1_624/A gnd INVX1_328/Y vdd INVX1
XOAI21X1_26 INVX1_27/A INVX1_29/Y INVX1_28/Y gnd OAI21X1_26/Y vdd OAI21X1
XAOI22X1_55 AOI22X1_55/A AND2X2_52/Y AOI22X1_55/C NOR2X1_71/Y gnd AOI22X1_55/Y vdd
+ AOI22X1
XNAND2X1_41 OAI21X1_23/Y AOI22X1_5/Y gnd NAND2X1_41/Y vdd NAND2X1
XAOI22X1_112 INVX1_378/A INVX1_377/Y INVX1_379/Y AOI22X1_112/D gnd OAI21X1_346/B vdd
+ AOI22X1
XDFFPOSX1_110 AOI22X1_55/C CLKBUF1_47/Y OAI21X1_166/Y gnd vdd DFFPOSX1
XINVX1_292 BUFX2_33/Y gnd INVX1_292/Y vdd INVX1
XDFFPOSX1_44 INVX1_58/A CLKBUF1_11/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XOAI21X1_471 INVX1_525/Y OAI21X1_471/B NOR2X1_203/Y gnd AOI21X1_76/C vdd OAI21X1
XAOI22X1_19 AOI22X1_19/A AND2X2_31/Y AOI22X1_19/C NOR2X1_32/Y gnd AOI22X1_19/Y vdd
+ AOI22X1
XOAI21X1_435 INVX1_483/Y OAI21X1_435/B NOR2X1_185/Y gnd AOI21X1_70/C vdd OAI21X1
XINVX1_256 INVX1_437/A gnd INVX1_256/Y vdd INVX1
XNAND3X1_82 BUFX2_51/Y INVX1_260/Y INVX1_261/Y gnd NAND3X1_82/Y vdd NAND3X1
XOAI21X1_399 INVX1_441/Y NAND2X1_386/Y NOR2X1_167/Y gnd AOI21X1_64/C vdd OAI21X1
XINVX1_220 AND2X2_59/B gnd INVX1_220/Y vdd INVX1
XNAND2X1_513 BUFX2_11/Y INVX1_601/Y gnd NAND2X1_513/Y vdd NAND2X1
XNAND3X1_46 BUFX2_50/Y NOR2X1_58/B INVX1_135/Y gnd NAND3X1_47/B vdd NAND3X1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XOAI21X1_363 INVX1_399/Y OAI21X1_363/B NOR2X1_149/Y gnd AOI21X1_58/C vdd OAI21X1
XCLKBUF1_5 BUFX2_4/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XNAND2X1_477 INVX1_553/A INVX1_554/A gnd NAND2X1_478/B vdd NAND2X1
XAND2X2_115 INVX1_522/A INVX1_508/A gnd AND2X2_115/Y vdd AND2X2
XNAND3X1_10 INVX1_5/A INVX1_39/A NAND3X1_8/C gnd OAI21X1_6/C vdd NAND3X1
XAND2X2_88 AND2X2_88/A AND2X2_88/B gnd AND2X2_88/Y vdd AND2X2
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_148 BUFX2_47/Y gnd NOR2X1_62/B vdd INVX1
XOAI21X1_327 INVX1_357/Y OAI21X1_327/B NOR2X1_131/Y gnd AOI21X1_52/C vdd OAI21X1
XNAND2X1_441 BUFX2_90/Y INVX1_513/A gnd OAI21X1_458/B vdd NAND2X1
XAND2X2_52 BUFX2_54/Y INVX1_178/A gnd AND2X2_52/Y vdd AND2X2
XFILL_23_1 gnd vdd FILL
XINVX1_112 AND2X2_4/B gnd INVX1_112/Y vdd INVX1
XFILL_14_1_1 gnd vdd FILL
XOAI21X1_291 INVX1_315/Y NAND2X1_287/Y NAND3X1_99/A gnd AOI21X1_46/C vdd OAI21X1
XNAND2X1_405 BUFX2_83/Y INVX1_464/Y gnd AOI22X1_136/D vdd NAND2X1
XFILL_12_3_2 gnd vdd FILL
XAND2X2_16 AND2X2_16/A NOR2X1_53/A gnd AND2X2_42/A vdd AND2X2
XNOR2X1_91 gnd INVX1_243/Y gnd NOR2X1_91/Y vdd NOR2X1
XOAI21X1_255 INVX1_277/Y AOI22X1_82/Y AOI22X1_83/Y gnd OAI21X1_255/Y vdd OAI21X1
XNAND2X1_369 INVX1_455/A INVX1_448/A gnd NOR3X1_4/C vdd NAND2X1
XINVX1_617 INVX1_160/A gnd INVX1_617/Y vdd INVX1
XNOR2X1_55 gnd NOR2X1_55/B gnd NOR2X1_55/Y vdd NOR2X1
XOAI21X1_219 INVX1_237/A INVX1_239/Y INVX1_238/Y gnd OAI21X1_220/C vdd OAI21X1
XNAND2X1_333 AND2X2_3/A NAND2X1_332/Y gnd NAND2X1_333/Y vdd NAND2X1
XCLKBUF1_43 BUFX2_1/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XINVX1_581 INVX1_581/A gnd INVX1_581/Y vdd INVX1
XNAND3X1_165 NOR2X1_215/Y NAND3X1_164/Y NAND3X1_165/C gnd NAND3X1_165/Y vdd NAND3X1
XNOR2X1_19 INVX1_16/A INVX1_17/Y gnd AOI22X1_4/B vdd NOR2X1
XOAI21X1_183 INVX1_197/A INVX1_195/Y OAI21X1_182/Y gnd NAND3X1_65/C vdd OAI21X1
XNOR2X1_216 NAND2X1_4/A INVX1_547/Y gnd NOR2X1_216/Y vdd NOR2X1
XNAND2X1_297 BUFX2_20/Y INVX1_328/Y gnd NAND2X1_297/Y vdd NAND2X1
XDFFPOSX1_363 AND2X2_49/B CLKBUF1_30/Y OAI21X1_550/Y gnd vdd DFFPOSX1
XFILL_3_0_0 gnd vdd FILL
XNAND3X1_129 NOR2X1_161/Y NAND3X1_128/Y OAI21X1_378/Y gnd NAND3X1_129/Y vdd NAND3X1
XBUFX2_130 NOR3X1_5/Y gnd BUFX2_130/Y vdd BUFX2
XINVX1_545 BUFX2_74/Y gnd INVX1_545/Y vdd INVX1
XFILL_21_1_1 gnd vdd FILL
XFILL_19_3_2 gnd vdd FILL
XOAI21X1_147 INVX1_153/Y INVX1_156/Y AOI22X1_49/C gnd OAI21X1_147/Y vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XNOR2X1_180 NAND2X1_8/A INVX1_463/Y gnd NOR2X1_180/Y vdd NOR2X1
XFILL_10_3 gnd vdd FILL
XNAND2X1_261 INVX1_282/A NAND2X1_261/B gnd AOI22X1_85/A vdd NAND2X1
XDFFPOSX1_327 INVX1_557/A CLKBUF1_47/Y OAI21X1_496/Y gnd vdd DFFPOSX1
XINVX1_509 BUFX2_30/Y gnd INVX1_509/Y vdd INVX1
XXNOR2X1_54 AND2X2_5/Y BUFX2_39/Y gnd AOI21X1_59/B vdd XNOR2X1
XOAI21X1_111 INVX1_115/Y NAND2X1_121/Y OAI21X1_111/C gnd DFFPOSX1_74/D vdd OAI21X1
XNOR2X1_144 INVX1_378/A INVX1_379/Y gnd NOR2X1_144/Y vdd NOR2X1
XNAND2X1_225 INVX1_237/A INVX1_240/Y gnd AOI22X1_72/D vdd NAND2X1
XDFFPOSX1_291 INVX1_241/A CLKBUF1_4/Y OAI21X1_442/Y gnd vdd DFFPOSX1
XINVX1_473 INVX1_473/A gnd INVX1_473/Y vdd INVX1
XXNOR2X1_18 BUFX2_47/Y AND2X2_7/Y gnd AOI21X1_23/B vdd XNOR2X1
XNAND2X1_189 AND2X2_8/Y INVX1_198/A gnd OAI21X1_185/B vdd NAND2X1
XNOR2X1_108 INVX1_294/A INVX1_295/Y gnd AOI22X1_89/D vdd NOR2X1
XDFFPOSX1_255 INVX1_431/A CLKBUF1_36/Y OAI21X1_388/Y gnd vdd DFFPOSX1
XAOI21X1_87 INVX1_604/Y XNOR2X1_82/Y AOI21X1_87/C gnd AOI21X1_87/Y vdd AOI21X1
XINVX1_437 INVX1_437/A gnd INVX1_437/Y vdd INVX1
XFILL_28_1_1 gnd vdd FILL
XBUFX2_90 BUFX2_88/A gnd BUFX2_90/Y vdd BUFX2
XNAND2X1_153 AND2X2_5/B BUFX2_47/Y gnd NAND2X1_153/Y vdd NAND2X1
XFILL_8_2_1 gnd vdd FILL
XFILL_26_3_2 gnd vdd FILL
XDFFPOSX1_219 INVX1_368/A CLKBUF1_43/Y OAI21X1_334/Y gnd vdd DFFPOSX1
XAOI21X1_51 INVX1_352/Y AOI21X1_51/B AOI21X1_51/C gnd AOI21X1_51/Y vdd AOI21X1
XINVX1_401 AND2X2_4/A gnd INVX1_401/Y vdd INVX1
XOAI21X1_4 INVX1_10/Y NOR3X1_1/Y OAI21X1_4/C gnd INVX1_178/A vdd OAI21X1
XBUFX2_54 BUFX2_54/A gnd BUFX2_54/Y vdd BUFX2
XNAND2X1_117 INVX1_106/A INVX1_104/Y gnd OAI21X1_106/B vdd NAND2X1
XOAI21X1_99 INVX1_98/Y OAI21X1_99/B NOR2X1_46/Y gnd OAI21X1_99/Y vdd OAI21X1
XINVX1_365 AND2X2_2/Y gnd INVX1_365/Y vdd INVX1
XAOI21X1_15 INVX1_100/Y XNOR2X1_10/Y OAI21X1_99/Y gnd AOI21X1_15/Y vdd AOI21X1
XOAI21X1_544 INVX1_613/Y AOI22X1_178/Y AOI22X1_179/Y gnd OAI21X1_544/Y vdd OAI21X1
XDFFPOSX1_183 AND2X2_72/B CLKBUF1_11/Y OAI21X1_279/Y gnd vdd DFFPOSX1
XBUFX2_18 BUFX2_18/A gnd BUFX2_18/Y vdd BUFX2
XNAND2X1_78 INVX1_56/A BUFX2_70/Y gnd NAND2X1_78/Y vdd NAND2X1
XAOI22X1_92 INVX1_308/A INVX1_307/Y INVX1_309/Y AOI22X1_92/D gnd AOI22X1_92/Y vdd
+ AOI22X1
XDFFPOSX1_147 INVX1_242/A CLKBUF1_31/Y OAI21X1_224/Y gnd vdd DFFPOSX1
XDFFPOSX1_81 NOR2X1_53/A CLKBUF1_1/Y NAND3X1_43/Y gnd vdd DFFPOSX1
XAOI22X1_149 AOI22X1_149/A AND2X2_117/Y AOI22X1_149/C NOR2X1_198/Y gnd AOI22X1_149/Y
+ vdd AOI22X1
XOAI21X1_63 INVX1_60/Y OAI21X1_63/B AOI22X1_21/Y gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_508 INVX1_571/Y OAI21X1_508/B OAI21X1_508/C gnd OAI21X1_508/Y vdd OAI21X1
XINVX1_329 AND2X2_21/B gnd INVX1_329/Y vdd INVX1
XAOI22X1_56 NOR2X1_73/A INVX1_181/Y NOR2X1_73/B AOI22X1_56/D gnd AOI22X1_56/Y vdd
+ AOI22X1
XOAI21X1_27 EN_response_get INVX1_27/Y OAI21X1_26/Y gnd OAI21X1_27/Y vdd OAI21X1
XNAND2X1_42 NAND2X1_42/A AOI22X1_6/Y gnd NAND2X1_42/Y vdd NAND2X1
XDFFPOSX1_45 INVX1_56/A CLKBUF1_11/Y NAND3X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 INVX1_171/A CLKBUF1_47/Y OAI21X1_168/Y gnd vdd DFFPOSX1
XAOI22X1_113 NAND2X1_341/Y AND2X2_90/Y AOI22X1_113/C NOR2X1_144/Y gnd OAI21X1_346/C
+ vdd AOI22X1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XOAI21X1_472 INVX1_529/Y AOI22X1_154/Y AOI22X1_155/Y gnd OAI21X1_472/Y vdd OAI21X1
XAOI22X1_20 INVX1_56/A INVX1_55/Y INVX1_57/Y AOI22X1_20/D gnd OAI21X1_63/B vdd AOI22X1
XOAI21X1_436 INVX1_487/Y AOI22X1_142/Y AOI22X1_143/Y gnd OAI21X1_436/Y vdd OAI21X1
XINVX1_257 BUFX2_33/Y gnd NOR2X1_96/B vdd INVX1
XNAND3X1_83 NOR2X1_96/Y NAND3X1_82/Y NAND3X1_83/C gnd NAND3X1_83/Y vdd NAND3X1
XOAI21X1_400 INVX1_445/Y OAI21X1_400/B OAI21X1_400/C gnd OAI21X1_400/Y vdd OAI21X1
XNAND2X1_514 INVX1_601/A INVX1_604/Y gnd AOI22X1_176/D vdd NAND2X1
XNAND3X1_47 NOR2X1_57/Y NAND3X1_47/B NAND3X1_47/C gnd NAND3X1_47/Y vdd NAND3X1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XINVX1_185 AND2X2_53/B gnd INVX1_185/Y vdd INVX1
XCLKBUF1_6 BUFX2_5/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XOAI21X1_364 INVX1_403/Y AOI22X1_118/Y AOI22X1_119/Y gnd OAI21X1_364/Y vdd OAI21X1
XAND2X2_116 INVX1_515/A INVX1_508/A gnd NOR2X1_196/B vdd AND2X2
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XNAND2X1_478 INVX1_555/A NAND2X1_478/B gnd AOI22X1_163/A vdd NAND2X1
XNAND3X1_11 INVX1_5/A INVX1_38/A NAND3X1_8/C gnd OAI21X1_7/C vdd NAND3X1
XAND2X2_89 AND2X2_87/B AND2X2_88/B gnd AND2X2_89/Y vdd AND2X2
XINVX1_31 OR2X2_2/B gnd INVX1_31/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XOAI21X1_328 INVX1_361/Y AOI22X1_106/Y AOI22X1_107/Y gnd OAI21X1_328/Y vdd OAI21X1
XNAND2X1_442 BUFX2_63/Y INVX1_510/Y gnd OAI21X1_459/B vdd NAND2X1
XAND2X2_53 INVX1_190/A AND2X2_53/B gnd AND2X2_53/Y vdd AND2X2
XFILL_23_2 gnd vdd FILL
XINVX1_113 INVX1_113/A gnd NOR2X1_51/B vdd INVX1
XOAI21X1_292 INVX1_319/Y AOI22X1_94/Y AOI22X1_95/Y gnd OAI21X1_292/Y vdd OAI21X1
XNAND2X1_406 NAND2X1_8/A INVX1_463/A gnd NAND2X1_406/Y vdd NAND2X1
XFILL_14_1_2 gnd vdd FILL
XAND2X2_17 INVX1_576/A AND2X2_17/B gnd INVX1_575/A vdd AND2X2
XNOR2X1_92 INVX1_245/A NOR2X1_92/B gnd NOR2X1_92/Y vdd NOR2X1
XOAI21X1_256 INVX1_279/A INVX1_281/Y INVX1_280/Y gnd OAI21X1_257/C vdd OAI21X1
XNAND2X1_370 BUFX2_80/Y INVX1_422/A gnd OAI21X1_380/B vdd NAND2X1
XINVX1_618 AND2X2_20/A gnd INVX1_618/Y vdd INVX1
XNOR2X1_56 NOR2X1_56/A NOR2X1_56/B gnd NOR2X1_56/Y vdd NOR2X1
XOAI21X1_220 BUFX2_17/Y INVX1_237/Y OAI21X1_220/C gnd NAND3X1_77/C vdd OAI21X1
XNAND2X1_334 INVX1_387/A INVX1_380/A gnd NOR3X1_3/A vdd NAND2X1
XFILL_15_2_0 gnd vdd FILL
XNAND3X1_166 BUFX2_94/Y INVX1_554/Y INVX1_555/Y gnd NAND3X1_166/Y vdd NAND3X1
XCLKBUF1_44 BUFX2_7/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XINVX1_582 INVX1_582/A gnd INVX1_582/Y vdd INVX1
XOAI21X1_184 INVX1_195/Y INVX1_198/Y AOI22X1_61/C gnd OAI21X1_185/C vdd OAI21X1
XNOR2X1_20 gnd INVX1_26/Y gnd NOR2X1_20/Y vdd NOR2X1
XNOR2X1_217 gnd INVX1_551/Y gnd NOR2X1_217/Y vdd NOR2X1
XNAND2X1_298 INVX1_624/A INVX1_331/Y gnd AOI22X1_98/D vdd NAND2X1
XDFFPOSX1_364 AND2X2_20/A CLKBUF1_50/Y AOI21X1_89/Y gnd vdd DFFPOSX1
XFILL_3_0_1 gnd vdd FILL
XNAND3X1_130 BUFX2_87/Y INVX1_428/Y INVX1_429/Y gnd NAND3X1_130/Y vdd NAND3X1
XBUFX2_131 NOR3X1_5/Y gnd INVX1_463/A vdd BUFX2
XINVX1_546 NAND2X1_4/A gnd INVX1_546/Y vdd INVX1
XFILL_21_1_2 gnd vdd FILL
XOAI21X1_148 INVX1_157/Y OAI21X1_148/B OAI21X1_147/Y gnd OAI21X1_148/Y vdd OAI21X1
XFILL_1_2_2 gnd vdd FILL
XNOR2X1_181 gnd INVX1_467/Y gnd NOR2X1_181/Y vdd NOR2X1
XNAND2X1_262 INVX1_575/A INVX1_289/A gnd OAI21X1_265/B vdd NAND2X1
XDFFPOSX1_328 INVX1_555/A CLKBUF1_47/Y AOI21X1_80/Y gnd vdd DFFPOSX1
XINVX1_510 BUFX2_89/Y gnd INVX1_510/Y vdd INVX1
XXNOR2X1_55 AND2X2_6/Y BUFX2_40/Y gnd AOI21X1_60/B vdd XNOR2X1
XNAND2X1_226 NOR2X1_90/A BUFX2_17/Y gnd NAND2X1_227/B vdd NAND2X1
XOAI21X1_112 INVX1_112/Y OAI21X1_112/B NOR2X1_50/Y gnd AOI21X1_17/C vdd OAI21X1
XNOR2X1_145 gnd INVX1_383/Y gnd NOR2X1_145/Y vdd NOR2X1
XDFFPOSX1_292 AND2X2_11/A CLKBUF1_17/Y AOI21X1_71/Y gnd vdd DFFPOSX1
XINVX1_474 BUFX2_34/Y gnd INVX1_474/Y vdd INVX1
XXNOR2X1_19 BUFX2_48/Y INVX1_160/A gnd XNOR2X1_19/Y vdd XNOR2X1
XFILL_22_2_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XNAND2X1_190 INVX1_197/A INVX1_195/Y gnd OAI21X1_186/B vdd NAND2X1
XNOR2X1_109 gnd INVX1_299/Y gnd NAND3X1_95/A vdd NOR2X1
XDFFPOSX1_256 INVX1_429/A CLKBUF1_10/Y AOI21X1_62/Y gnd vdd DFFPOSX1
XAOI21X1_88 INVX1_611/Y AOI21X1_88/B AOI21X1_88/C gnd AOI21X1_88/Y vdd AOI21X1
XINVX1_438 AND2X2_96/A gnd INVX1_438/Y vdd INVX1
XFILL_28_1_2 gnd vdd FILL
XBUFX2_91 BUFX2_88/A gnd BUFX2_91/Y vdd BUFX2
XNAND2X1_154 INVX1_149/A NAND2X1_153/Y gnd AOI22X1_47/A vdd NAND2X1
XFILL_8_2_2 gnd vdd FILL
XDFFPOSX1_220 AND2X2_2/A CLKBUF1_30/Y AOI21X1_53/Y gnd vdd DFFPOSX1
XINVX1_402 INVX1_402/A gnd INVX1_402/Y vdd INVX1
XAOI21X1_52 INVX1_359/Y AOI21X1_52/B AOI21X1_52/C gnd AOI21X1_52/Y vdd AOI21X1
XBUFX2_55 BUFX2_54/A gnd BUFX2_55/Y vdd BUFX2
XNAND2X1_118 AND2X2_2/Y INVX1_107/Y gnd AOI22X1_34/D vdd NAND2X1
XOAI21X1_5 INVX1_11/Y NOR3X1_1/Y NAND3X1_9/Y gnd AND2X2_59/B vdd OAI21X1
XDFFPOSX1_184 AND2X2_71/B CLKBUF1_38/Y AOI21X1_44/Y gnd vdd DFFPOSX1
XAOI21X1_16 INVX1_107/Y AOI21X1_16/B AOI21X1_16/C gnd AOI21X1_16/Y vdd AOI21X1
XINVX1_366 AND2X2_2/A gnd INVX1_366/Y vdd INVX1
XOAI21X1_545 BUFX2_8/Y INVX1_617/Y INVX1_616/Y gnd OAI21X1_546/C vdd OAI21X1
XFILL_14_1 gnd vdd FILL
XBUFX2_19 BUFX2_18/A gnd BUFX2_19/Y vdd BUFX2
XOAI21X1_64 INVX1_67/A INVX1_81/A INVX1_74/A gnd NAND2X1_81/B vdd OAI21X1
XNAND2X1_79 INVX1_58/A NAND2X1_78/Y gnd NAND2X1_79/Y vdd NAND2X1
XAOI22X1_93 AOI22X1_93/A AND2X2_74/Y AOI22X1_93/C NOR2X1_112/Y gnd AOI22X1_93/Y vdd
+ AOI22X1
XDFFPOSX1_148 INVX1_240/A CLKBUF1_16/Y AOI21X1_35/Y gnd vdd DFFPOSX1
XFILL_9_3_0 gnd vdd FILL
XDFFPOSX1_82 AOI22X1_41/C CLKBUF1_50/Y DFFPOSX1_82/D gnd vdd DFFPOSX1
XAOI22X1_150 INVX1_511/A INVX1_510/Y INVX1_512/Y NAND2X1_443/Y gnd OAI21X1_460/B vdd
+ AOI22X1
XINVX1_330 BUFX2_20/Y gnd INVX1_330/Y vdd INVX1
XOAI21X1_509 BUFX2_124/Y INVX1_575/Y INVX1_574/Y gnd OAI21X1_510/C vdd OAI21X1
XAOI22X1_57 AOI22X1_57/A AND2X2_53/Y AOI22X1_57/C NOR2X1_73/Y gnd AOI22X1_57/Y vdd
+ AOI22X1
XOAI21X1_28 INVX1_30/Y NOR2X1_21/Y NAND2X1_45/Y gnd OAI21X1_28/Y vdd OAI21X1
XNAND2X1_43 NAND2X1_43/A AOI22X1_7/Y gnd NAND2X1_43/Y vdd NAND2X1
XDFFPOSX1_46 OAI21X1_67/C CLKBUF1_25/Y OAI21X1_68/Y gnd vdd DFFPOSX1
XAOI22X1_114 INVX1_385/A INVX1_384/Y INVX1_386/Y AOI22X1_114/D gnd OAI21X1_352/B vdd
+ AOI22X1
XINVX1_294 INVX1_294/A gnd INVX1_294/Y vdd INVX1
XDFFPOSX1_112 AND2X2_50/B CLKBUF1_32/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XOAI21X1_473 BUFX2_62/Y INVX1_533/Y INVX1_532/Y gnd OAI21X1_473/Y vdd OAI21X1
XAOI22X1_21 NAND2X1_79/Y AND2X2_32/Y AOI22X1_21/C NOR2X1_34/Y gnd AOI22X1_21/Y vdd
+ AOI22X1
XDFFPOSX1_10 INVX1_25/A CLKBUF1_18/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XOAI21X1_437 BUFX2_129/Y INVX1_491/Y INVX1_490/Y gnd OAI21X1_437/Y vdd OAI21X1
XINVX1_258 BUFX2_51/Y gnd INVX1_258/Y vdd INVX1
XNAND3X1_84 BUFX2_60/Y NOR2X1_99/B INVX1_268/Y gnd NAND3X1_84/Y vdd NAND3X1
XINVX1_222 BUFX2_31/Y gnd INVX1_222/Y vdd INVX1
XOAI21X1_401 BUFX2_113/Y INVX1_449/Y INVX1_448/Y gnd OAI21X1_402/C vdd OAI21X1
XNAND3X1_48 BUFX2_46/Y INVX1_141/Y INVX1_142/Y gnd NAND3X1_48/Y vdd NAND3X1
XNAND2X1_515 INVX1_602/A BUFX2_11/Y gnd NAND2X1_516/B vdd NAND2X1
XINVX1_68 BUFX2_32/Y gnd INVX1_68/Y vdd INVX1
XOAI21X1_365 BUFX2_39/Y INVX1_407/Y INVX1_406/Y gnd OAI21X1_365/Y vdd OAI21X1
XINVX1_186 OR2X2_4/A gnd INVX1_186/Y vdd INVX1
XAND2X2_117 BUFX2_25/Y INVX1_46/A gnd AND2X2_117/Y vdd AND2X2
XCLKBUF1_7 BUFX2_7/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XNAND2X1_479 BUFX2_99/Y INVX1_562/A gnd NAND2X1_479/Y vdd NAND2X1
XNAND3X1_12 BUFX2_30/Y NAND2X1_26/Y NAND3X1_12/C gnd DFFPOSX1_1/D vdd NAND3X1
XAND2X2_90 BUFX2_73/Y INVX1_88/A gnd AND2X2_90/Y vdd AND2X2
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XFILL_10_0_0 gnd vdd FILL
XFILL_1_2 gnd vdd FILL
XINVX1_150 AND2X2_47/B gnd INVX1_150/Y vdd INVX1
XOAI21X1_329 INVX1_363/A INVX1_365/Y INVX1_364/Y gnd OAI21X1_330/C vdd OAI21X1
XNAND2X1_443 BUFX2_89/Y INVX1_513/Y gnd NAND2X1_443/Y vdd NAND2X1
XAND2X2_54 AND2X2_3/Y INVX1_375/A gnd AND2X2_54/Y vdd AND2X2
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XOAI21X1_293 INVX1_582/A INVX1_323/Y INVX1_322/Y gnd OAI21X1_293/Y vdd OAI21X1
XNAND2X1_407 INVX1_464/A NAND2X1_406/Y gnd AOI22X1_137/A vdd NAND2X1
XAND2X2_18 INVX1_583/A AND2X2_18/B gnd INVX1_582/A vdd AND2X2
XNOR2X1_93 NOR2X1_93/A NOR2X1_93/B gnd BUFX2_58/A vdd NOR2X1
XOAI21X1_257 BUFX2_59/Y INVX1_279/Y OAI21X1_257/C gnd NAND3X1_89/C vdd OAI21X1
XNAND2X1_371 INVX1_421/A INVX1_419/Y gnd OAI21X1_381/B vdd NAND2X1
XINVX1_619 INVX1_619/A gnd INVX1_619/Y vdd INVX1
XNOR2X1_57 gnd NOR2X1_57/B gnd NOR2X1_57/Y vdd NOR2X1
XOAI21X1_221 INVX1_237/Y INVX1_240/Y AOI22X1_73/C gnd OAI21X1_222/C vdd OAI21X1
XNAND2X1_335 INVX1_399/A INVX1_394/A gnd NOR3X1_3/B vdd NAND2X1
XFILL_15_2_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XCLKBUF1_45 BUFX2_5/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XNAND3X1_167 NOR2X1_217/Y NAND3X1_166/Y OAI21X1_492/Y gnd NAND3X1_167/Y vdd NAND3X1
XINVX1_583 INVX1_583/A gnd INVX1_583/Y vdd INVX1
XOAI21X1_185 INVX1_199/Y OAI21X1_185/B OAI21X1_185/C gnd OAI21X1_185/Y vdd OAI21X1
XNOR2X1_21 INVX1_27/Y INVX1_31/Y gnd NOR2X1_21/Y vdd NOR2X1
XNOR2X1_218 INVX1_553/A INVX1_554/Y gnd NOR2X1_218/Y vdd NOR2X1
XNAND2X1_299 AND2X2_21/B BUFX2_20/Y gnd NAND2X1_300/B vdd NAND2X1
XNAND3X1_131 NOR2X1_163/Y NAND3X1_130/Y OAI21X1_384/Y gnd NAND3X1_131/Y vdd NAND3X1
XDFFPOSX1_365 INVX1_616/A CLKBUF1_50/Y NAND3X1_185/Y gnd vdd DFFPOSX1
XINVX1_547 INVX1_547/A gnd INVX1_547/Y vdd INVX1
XFILL_3_0_2 gnd vdd FILL
XBUFX2_132 NOR3X1_5/Y gnd BUFX2_132/Y vdd BUFX2
XOAI21X1_149 INVX1_154/Y OAI21X1_149/B NOR2X1_63/Y gnd AOI21X1_23/C vdd OAI21X1
XNOR2X1_182 INVX1_469/A INVX1_470/Y gnd NOR2X1_182/Y vdd NOR2X1
XNAND2X1_263 BUFX2_57/Y INVX1_286/Y gnd NAND2X1_263/Y vdd NAND2X1
XDFFPOSX1_329 INVX1_553/A CLKBUF1_29/Y NAND3X1_167/Y gnd vdd DFFPOSX1
XINVX1_511 INVX1_511/A gnd INVX1_511/Y vdd INVX1
XOAI21X1_113 INVX1_116/Y AOI22X1_36/Y AOI22X1_37/Y gnd OAI21X1_113/Y vdd OAI21X1
XXNOR2X1_56 INVX1_421/A BUFX2_79/Y gnd XNOR2X1_56/Y vdd XNOR2X1
XNAND2X1_227 INVX1_240/A NAND2X1_227/B gnd AOI22X1_73/A vdd NAND2X1
XNOR2X1_146 INVX1_385/A INVX1_386/Y gnd NOR2X1_146/Y vdd NOR2X1
XDFFPOSX1_293 INVX1_490/A CLKBUF1_31/Y NAND3X1_149/Y gnd vdd DFFPOSX1
XINVX1_475 INVX1_475/A gnd INVX1_475/Y vdd INVX1
XFILL_24_0_0 gnd vdd FILL
XXNOR2X1_20 BUFX2_85/Y INVX1_167/A gnd AOI21X1_25/B vdd XNOR2X1
XFILL_4_1_0 gnd vdd FILL
XFILL_22_2_1 gnd vdd FILL
XNOR2X1_110 INVX1_301/A INVX1_302/Y gnd AOI22X1_91/D vdd NOR2X1
XNAND2X1_191 AND2X2_8/Y INVX1_198/Y gnd AOI22X1_60/D vdd NAND2X1
XFILL_2_3_1 gnd vdd FILL
XINVX1_439 BUFX2_28/Y gnd INVX1_439/Y vdd INVX1
XDFFPOSX1_257 INVX1_427/A CLKBUF1_33/Y NAND3X1_131/Y gnd vdd DFFPOSX1
XAOI21X1_89 INVX1_618/Y XNOR2X1_84/Y AOI21X1_89/C gnd AOI21X1_89/Y vdd AOI21X1
XBUFX2_92 BUFX2_88/A gnd BUFX2_92/Y vdd BUFX2
XNAND2X1_155 AND2X2_7/Y INVX1_156/A gnd OAI21X1_148/B vdd NAND2X1
XAOI21X1_53 INVX1_366/Y AOI21X1_53/B AOI21X1_53/C gnd AOI21X1_53/Y vdd AOI21X1
XDFFPOSX1_221 INVX1_364/A CLKBUF1_30/Y NAND3X1_113/Y gnd vdd DFFPOSX1
XINVX1_403 INVX1_115/A gnd INVX1_403/Y vdd INVX1
XBUFX2_56 BUFX2_54/A gnd BUFX2_56/Y vdd BUFX2
XNAND2X1_119 AND2X2_2/B INVX1_106/A gnd NAND2X1_119/Y vdd NAND2X1
XOAI21X1_6 INVX1_12/Y NOR3X1_1/Y OAI21X1_6/C gnd AND2X2_66/B vdd OAI21X1
XAOI21X1_17 INVX1_114/Y AOI21X1_17/B AOI21X1_17/C gnd AOI21X1_17/Y vdd AOI21X1
XDFFPOSX1_185 INVX1_301/A CLKBUF1_38/Y NAND3X1_95/Y gnd vdd DFFPOSX1
XINVX1_367 INVX1_367/A gnd INVX1_367/Y vdd INVX1
XOAI21X1_546 INVX1_160/A INVX1_615/Y OAI21X1_546/C gnd OAI21X1_546/Y vdd OAI21X1
XFILL_14_2 gnd vdd FILL
XBUFX2_20 BUFX2_18/A gnd BUFX2_20/Y vdd BUFX2
XAOI22X1_94 AND2X2_12/B INVX1_314/Y INVX1_316/Y AOI22X1_94/D gnd AOI22X1_94/Y vdd
+ AOI22X1
XDFFPOSX1_83 AND2X2_99/B CLKBUF1_50/Y OAI21X1_125/Y gnd vdd DFFPOSX1
XNAND2X1_80 INVX1_67/A INVX1_81/A gnd NAND2X1_80/Y vdd NAND2X1
XOAI21X1_65 AND2X2_1/Y INVX1_64/Y INVX1_63/Y gnd OAI21X1_66/C vdd OAI21X1
XDFFPOSX1_149 NOR2X1_90/A CLKBUF1_31/Y NAND3X1_77/Y gnd vdd DFFPOSX1
XFILL_9_3_1 gnd vdd FILL
XAOI22X1_151 AOI22X1_151/A AND2X2_118/Y AOI22X1_151/C NOR2X1_200/Y gnd AOI22X1_151/Y
+ vdd AOI22X1
XOAI21X1_510 INVX1_575/A INVX1_573/Y OAI21X1_510/C gnd NAND3X1_173/C vdd OAI21X1
XINVX1_331 INVX1_331/A gnd INVX1_331/Y vdd INVX1
XAOI22X1_58 AND2X2_3/B INVX1_188/Y NOR2X1_75/B AOI22X1_58/D gnd AOI22X1_58/Y vdd AOI22X1
XOAI21X1_29 INVX1_32/Y NOR2X1_21/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XNAND2X1_44 INVX1_27/A INVX1_29/Y gnd OR2X2_2/A vdd NAND2X1
XDFFPOSX1_47 INVX1_67/A CLKBUF1_26/Y OAI21X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 NOR2X1_71/A CLKBUF1_9/Y NAND3X1_59/Y gnd vdd DFFPOSX1
XAOI22X1_115 AOI22X1_115/A AND2X2_91/Y OAI21X1_349/C NOR2X1_146/Y gnd AOI22X1_115/Y
+ vdd AOI22X1
XINVX1_295 BUFX2_100/Y gnd INVX1_295/Y vdd INVX1
XOAI21X1_474 INVX1_244/A INVX1_531/Y OAI21X1_473/Y gnd OAI21X1_474/Y vdd OAI21X1
XAOI22X1_22 AND2X2_1/B INVX1_62/Y INVX1_64/Y NAND2X1_84/Y gnd AOI22X1_22/Y vdd AOI22X1
XDFFPOSX1_11 INVX1_6/A CLKBUF1_18/Y NAND2X1_37/Y gnd vdd DFFPOSX1
XINVX1_259 NOR2X1_97/A gnd INVX1_259/Y vdd INVX1
XOAI21X1_438 INVX1_237/A INVX1_489/Y OAI21X1_437/Y gnd OAI21X1_438/Y vdd OAI21X1
XNAND3X1_85 NOR2X1_98/Y NAND3X1_84/Y NAND3X1_85/C gnd NAND3X1_85/Y vdd NAND3X1
XINVX1_223 BUFX2_16/Y gnd INVX1_223/Y vdd INVX1
XOAI21X1_402 AND2X2_8/Y INVX1_447/Y OAI21X1_402/C gnd NAND3X1_137/C vdd OAI21X1
XNAND3X1_49 NOR2X1_59/Y NAND3X1_48/Y NAND3X1_49/C gnd NAND3X1_49/Y vdd NAND3X1
XNAND2X1_516 INVX1_604/A NAND2X1_516/B gnd AOI22X1_177/A vdd NAND2X1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XINVX1_187 BUFX2_31/Y gnd NOR2X1_74/B vdd INVX1
XOAI21X1_366 AND2X2_5/Y INVX1_405/Y OAI21X1_365/Y gnd OAI21X1_366/Y vdd OAI21X1
XCLKBUF1_8 BUFX2_1/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XAND2X2_118 BUFX2_90/Y INVX1_395/A gnd AND2X2_118/Y vdd AND2X2
XNAND2X1_480 BUFX2_125/Y INVX1_559/Y gnd OAI21X1_501/B vdd NAND2X1
XNAND3X1_13 NOR2X1_16/Y OAI21X1_9/Y OR2X2_1/Y gnd NAND3X1_13/Y vdd NAND3X1
XAND2X2_91 BUFX2_79/Y AND2X2_99/B gnd AND2X2_91/Y vdd AND2X2
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XOAI21X1_330 AND2X2_2/Y INVX1_363/Y OAI21X1_330/C gnd NAND3X1_113/C vdd OAI21X1
XFILL_10_0_1 gnd vdd FILL
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XNAND2X1_444 INVX1_511/A BUFX2_61/Y gnd NAND2X1_445/B vdd NAND2X1
XAND2X2_55 AND2X2_8/Y INVX1_199/A gnd AND2X2_55/Y vdd AND2X2
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XOAI21X1_294 BUFX2_19/Y INVX1_321/Y OAI21X1_293/Y gnd OAI21X1_294/Y vdd OAI21X1
XNAND2X1_408 BUFX2_91/Y INVX1_471/A gnd NAND2X1_408/Y vdd NAND2X1
XAND2X2_19 INVX1_611/A INVX1_77/A gnd INVX1_76/A vdd AND2X2
XNOR2X1_94 gnd INVX1_250/Y gnd NOR2X1_94/Y vdd NOR2X1
XOAI21X1_258 INVX1_279/Y INVX1_282/Y AOI22X1_85/C gnd OAI21X1_259/C vdd OAI21X1
XNAND2X1_372 BUFX2_80/Y INVX1_422/Y gnd AOI22X1_124/D vdd NAND2X1
XINVX1_620 AND2X2_49/B gnd INVX1_620/Y vdd INVX1
XOAI21X1_222 INVX1_241/Y OAI21X1_222/B OAI21X1_222/C gnd OAI21X1_222/Y vdd OAI21X1
XNOR2X1_58 INVX1_133/A NOR2X1_58/B gnd NOR2X1_58/Y vdd NOR2X1
XNAND2X1_336 INVX1_413/A INVX1_406/A gnd NOR3X1_3/C vdd NAND2X1
XFILL_17_0_1 gnd vdd FILL
XFILL_15_2_2 gnd vdd FILL
XNOR2X1_22 INVX1_27/A INVX1_28/Y gnd NOR2X1_22/Y vdd NOR2X1
XNAND3X1_168 BUFX2_99/Y INVX1_561/Y INVX1_562/Y gnd NAND3X1_169/B vdd NAND3X1
XINVX1_584 INVX1_584/A gnd INVX1_584/Y vdd INVX1
XCLKBUF1_46 BUFX2_6/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XOAI21X1_186 INVX1_196/Y OAI21X1_186/B NOR2X1_76/Y gnd AOI21X1_29/C vdd OAI21X1
XNOR2X1_219 gnd INVX1_558/Y gnd NOR2X1_219/Y vdd NOR2X1
XNAND2X1_300 INVX1_331/A NAND2X1_300/B gnd AOI22X1_99/A vdd NAND2X1
XCLKBUF1_10 BUFX2_1/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XBUFX2_133 NOR3X1_5/Y gnd BUFX2_133/Y vdd BUFX2
XNAND3X1_132 BUFX2_96/Y INVX1_435/Y INVX1_436/Y gnd NAND3X1_132/Y vdd NAND3X1
XINVX1_548 INVX1_548/A gnd INVX1_548/Y vdd INVX1
XDFFPOSX1_366 AOI22X1_183/C CLKBUF1_7/Y OAI21X1_554/Y gnd vdd DFFPOSX1
XOAI21X1_150 INVX1_158/Y AOI22X1_48/Y AOI22X1_49/Y gnd DFFPOSX1_99/D vdd OAI21X1
XNOR2X1_183 gnd INVX1_474/Y gnd NOR2X1_183/Y vdd NOR2X1
XNAND2X1_264 INVX1_575/A INVX1_289/Y gnd AOI22X1_86/D vdd NAND2X1
XDFFPOSX1_330 OAI21X1_499/C CLKBUF1_47/Y OAI21X1_500/Y gnd vdd DFFPOSX1
XFILL_27_1 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XINVX1_512 BUFX2_63/Y gnd INVX1_512/Y vdd INVX1
XXNOR2X1_57 BUFX2_116/Y BUFX2_87/Y gnd AOI21X1_62/B vdd XNOR2X1
XOAI21X1_114 AND2X2_42/A NOR2X1_53/B INVX1_119/Y gnd OAI21X1_115/C vdd OAI21X1
XNAND2X1_228 INVX1_244/A INVX1_247/A gnd NAND2X1_228/Y vdd NAND2X1
XNOR2X1_147 gnd INVX1_390/Y gnd NOR2X1_147/Y vdd NOR2X1
XDFFPOSX1_294 OAI21X1_445/C CLKBUF1_23/Y OAI21X1_446/Y gnd vdd DFFPOSX1
XINVX1_476 INVX1_476/A gnd INVX1_476/Y vdd INVX1
XFILL_24_0_1 gnd vdd FILL
XFILL_22_2_2 gnd vdd FILL
XFILL_2_3_2 gnd vdd FILL
XFILL_4_1_1 gnd vdd FILL
XXNOR2X1_21 INVX1_167/A BUFX2_54/Y gnd AOI21X1_26/B vdd XNOR2X1
XNOR2X1_111 gnd INVX1_306/Y gnd NOR2X1_111/Y vdd NOR2X1
XNAND2X1_192 AND2X2_8/B INVX1_197/A gnd NAND2X1_193/B vdd NAND2X1
XINVX1_440 INVX1_440/A gnd INVX1_440/Y vdd INVX1
XDFFPOSX1_258 AOI22X1_129/C CLKBUF1_17/Y OAI21X1_392/Y gnd vdd DFFPOSX1
XAOI21X1_90 INVX1_625/Y XNOR2X1_85/Y AOI21X1_90/C gnd AOI21X1_90/Y vdd AOI21X1
XBUFX2_93 BUFX2_96/A gnd BUFX2_93/Y vdd BUFX2
XNAND2X1_156 BUFX2_49/Y INVX1_153/Y gnd OAI21X1_149/B vdd NAND2X1
XAOI21X1_54 INVX1_373/Y XNOR2X1_49/Y AOI21X1_54/C gnd AOI21X1_54/Y vdd AOI21X1
XDFFPOSX1_222 OAI21X1_337/C CLKBUF1_10/Y OAI21X1_338/Y gnd vdd DFFPOSX1
XINVX1_404 BUFX2_35/Y gnd INVX1_404/Y vdd INVX1
XBUFX2_57 BUFX2_58/A gnd BUFX2_57/Y vdd BUFX2
XNAND2X1_120 INVX1_107/A NAND2X1_119/Y gnd AOI22X1_35/A vdd NAND2X1
XFILL_23_3_0 gnd vdd FILL
XOAI21X1_7 INVX1_13/Y NOR3X1_1/Y OAI21X1_7/C gnd AND2X2_73/B vdd OAI21X1
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XAOI21X1_18 INVX1_121/Y AOI21X1_18/B AOI21X1_18/C gnd AOI21X1_18/Y vdd AOI21X1
XDFFPOSX1_186 AOI22X1_93/C CLKBUF1_40/Y OAI21X1_283/Y gnd vdd DFFPOSX1
XOAI21X1_547 INVX1_615/Y INVX1_618/Y AOI22X1_181/C gnd OAI21X1_547/Y vdd OAI21X1
XBUFX2_21 BUFX2_18/A gnd BUFX2_21/Y vdd BUFX2
XAOI22X1_95 AOI22X1_95/A AND2X2_75/Y AOI22X1_95/C AOI22X1_95/D gnd AOI22X1_95/Y vdd
+ AOI22X1
XDFFPOSX1_84 NAND2X1_5/B CLKBUF1_50/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XNAND2X1_81 NAND2X1_80/Y NAND2X1_81/B gnd INVX1_59/A vdd NAND2X1
XOAI21X1_66 INVX1_64/A INVX1_62/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XFILL_9_3_2 gnd vdd FILL
XDFFPOSX1_150 AOI22X1_75/C CLKBUF1_35/Y OAI21X1_228/Y gnd vdd DFFPOSX1
XINVX1_332 INVX1_627/A gnd INVX1_332/Y vdd INVX1
XOAI21X1_511 INVX1_573/Y INVX1_576/Y AOI22X1_169/C gnd OAI21X1_512/C vdd OAI21X1
XAOI22X1_152 INVX1_518/A INVX1_517/Y INVX1_519/Y NAND2X1_448/Y gnd AOI22X1_152/Y vdd
+ AOI22X1
XAOI22X1_59 AOI22X1_59/A AND2X2_54/Y AOI22X1_59/C NOR2X1_75/Y gnd AOI22X1_59/Y vdd
+ AOI22X1
XNAND2X1_45 OR2X2_5/A NOR2X1_21/Y gnd NAND2X1_45/Y vdd NAND2X1
XDFFPOSX1_114 AOI22X1_57/C CLKBUF1_49/Y OAI21X1_172/Y gnd vdd DFFPOSX1
XOAI21X1_30 INVX1_33/Y NOR2X1_21/Y NAND2X1_47/Y gnd OAI21X1_30/Y vdd OAI21X1
XDFFPOSX1_48 INVX1_65/A CLKBUF1_26/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XAOI22X1_116 INVX1_392/A INVX1_391/Y INVX1_393/Y AOI22X1_116/D gnd OAI21X1_358/B vdd
+ AOI22X1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XOAI21X1_475 INVX1_531/Y INVX1_534/Y OAI21X1_475/C gnd OAI21X1_476/C vdd OAI21X1
XAOI22X1_23 AOI22X1_23/A AND2X2_33/Y OAI21X1_67/C NOR2X1_36/Y gnd AOI22X1_23/Y vdd
+ AOI22X1
XDFFPOSX1_12 INVX1_8/A CLKBUF1_34/Y NAND2X1_38/Y gnd vdd DFFPOSX1
XOAI21X1_439 INVX1_489/Y INVX1_492/Y AOI22X1_145/C gnd OAI21X1_440/C vdd OAI21X1
XINVX1_260 INVX1_251/A gnd INVX1_260/Y vdd INVX1
XNAND3X1_86 AND2X2_9/Y INVX1_274/Y INVX1_275/Y gnd NAND3X1_86/Y vdd NAND3X1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XOAI21X1_403 INVX1_447/Y INVX1_450/Y AOI22X1_133/C gnd OAI21X1_404/C vdd OAI21X1
XNAND3X1_50 AND2X2_5/Y NOR2X1_62/B INVX1_149/Y gnd NAND3X1_51/B vdd NAND3X1
XNAND2X1_517 BUFX2_9/Y INVX1_611/A gnd NAND2X1_517/Y vdd NAND2X1
XINVX1_188 AND2X2_3/Y gnd INVX1_188/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XOAI21X1_367 INVX1_405/Y INVX1_408/Y AOI22X1_121/C gnd OAI21X1_367/Y vdd OAI21X1
XNAND2X1_481 BUFX2_98/Y INVX1_562/Y gnd AOI22X1_164/D vdd NAND2X1
XAND2X2_119 BUFX2_94/Y INVX1_437/A gnd AND2X2_119/Y vdd AND2X2
XNAND3X1_14 INVX1_16/A INVX1_3/Y EN_request_put gnd OAI21X1_19/C vdd NAND3X1
XCLKBUF1_9 BUFX2_4/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XAND2X2_92 BUFX2_92/Y INVX1_395/A gnd AND2X2_92/Y vdd AND2X2
XINVX1_152 BUFX2_35/Y gnd INVX1_152/Y vdd INVX1
XOAI21X1_331 INVX1_363/Y INVX1_366/Y OAI21X1_331/C gnd OAI21X1_331/Y vdd OAI21X1
XFILL_10_0_2 gnd vdd FILL
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XNAND2X1_445 INVX1_513/A NAND2X1_445/B gnd AOI22X1_151/A vdd NAND2X1
XAND2X2_56 INVX1_484/A INVX1_487/A gnd AND2X2_56/Y vdd AND2X2
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XOAI21X1_295 INVX1_321/Y INVX1_324/Y AOI22X1_97/C gnd OAI21X1_296/C vdd OAI21X1
XNAND2X1_409 BUFX2_132/Y INVX1_468/Y gnd NAND2X1_409/Y vdd NAND2X1
XAND2X2_20 AND2X2_20/A INVX1_161/A gnd INVX1_160/A vdd AND2X2
XNOR2X1_95 NOR2X1_95/A INVX1_253/Y gnd NOR2X1_95/Y vdd NOR2X1
XOAI21X1_259 INVX1_283/Y NAND2X1_257/Y OAI21X1_259/C gnd OAI21X1_259/Y vdd OAI21X1
XNAND2X1_373 INVX1_420/A INVX1_421/A gnd NAND2X1_373/Y vdd NAND2X1
XFILL_11_1_0 gnd vdd FILL
XINVX1_621 INVX1_89/A gnd INVX1_621/Y vdd INVX1
XOAI21X1_223 INVX1_238/Y OAI21X1_223/B NOR2X1_89/Y gnd AOI21X1_35/C vdd OAI21X1
XNOR2X1_59 gnd NOR2X1_59/B gnd NOR2X1_59/Y vdd NOR2X1
XNAND2X1_337 BUFX2_73/Y INVX1_380/A gnd OAI21X1_344/B vdd NAND2X1
XFILL_17_0_2 gnd vdd FILL
XNAND3X1_169 NOR2X1_219/Y NAND3X1_169/B NAND3X1_169/C gnd NAND3X1_169/Y vdd NAND3X1
XINVX1_585 INVX1_325/A gnd INVX1_585/Y vdd INVX1
XNOR2X1_23 INVX1_28/A INVX1_29/Y gnd AOI22X1_9/B vdd NOR2X1
XCLKBUF1_47 BUFX2_2/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XOAI21X1_187 INVX1_200/Y AOI22X1_60/Y AOI22X1_61/Y gnd OAI21X1_187/Y vdd OAI21X1
XNOR2X1_220 INVX1_560/A INVX1_561/Y gnd NOR2X1_220/Y vdd NOR2X1
XNAND2X1_301 INVX1_345/A INVX1_338/A gnd NOR3X1_2/A vdd NAND2X1
XBUFX2_134 NOR3X1_5/Y gnd BUFX2_134/Y vdd BUFX2
XFILL_5_1 gnd vdd FILL
XNAND3X1_133 NOR2X1_165/Y NAND3X1_132/Y NAND3X1_133/C gnd NAND3X1_133/Y vdd NAND3X1
XINVX1_549 INVX1_88/A gnd INVX1_549/Y vdd INVX1
XDFFPOSX1_367 INVX1_627/A CLKBUF1_7/Y OAI21X1_556/Y gnd vdd DFFPOSX1
XCLKBUF1_11 BUFX2_6/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XOAI21X1_151 INVX1_160/A INVX1_162/Y INVX1_161/Y gnd OAI21X1_152/C vdd OAI21X1
XNOR2X1_184 INVX1_476/A INVX1_477/Y gnd NOR2X1_184/Y vdd NOR2X1
XNAND2X1_265 AND2X2_17/B BUFX2_57/Y gnd NAND2X1_265/Y vdd NAND2X1
XDFFPOSX1_331 INVX1_564/A CLKBUF1_42/Y OAI21X1_502/Y gnd vdd DFFPOSX1
XFILL_18_1_0 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XINVX1_513 INVX1_513/A gnd INVX1_513/Y vdd INVX1
XOAI21X1_115 BUFX2_105/Y INVX1_118/Y OAI21X1_115/C gnd NAND3X1_43/C vdd OAI21X1
XXNOR2X1_58 BUFX2_112/Y BUFX2_96/Y gnd XNOR2X1_58/Y vdd XNOR2X1
XNOR2X1_148 INVX1_392/A INVX1_393/Y gnd NOR2X1_148/Y vdd NOR2X1
XNAND2X1_229 BUFX2_15/Y INVX1_244/Y gnd OAI21X1_229/B vdd NAND2X1
XINVX1_477 BUFX2_133/Y gnd INVX1_477/Y vdd INVX1
XDFFPOSX1_295 INVX1_501/A CLKBUF1_19/Y OAI21X1_448/Y gnd vdd DFFPOSX1
XXNOR2X1_22 BUFX2_67/Y BUFX2_108/Y gnd AOI21X1_27/B vdd XNOR2X1
XFILL_24_0_2 gnd vdd FILL
XNAND2X1_193 INVX1_198/A NAND2X1_193/B gnd AOI22X1_61/A vdd NAND2X1
XFILL_4_1_2 gnd vdd FILL
XNOR2X1_112 INVX1_308/A INVX1_309/Y gnd NOR2X1_112/Y vdd NOR2X1
XDFFPOSX1_259 AND2X2_96/A CLKBUF1_35/Y OAI21X1_394/Y gnd vdd DFFPOSX1
XINVX1_441 INVX1_441/A gnd INVX1_441/Y vdd INVX1
XBUFX2_94 BUFX2_96/A gnd BUFX2_94/Y vdd BUFX2
XNAND2X1_157 AND2X2_7/Y INVX1_156/Y gnd AOI22X1_48/D vdd NAND2X1
XDFFPOSX1_223 INVX1_375/A CLKBUF1_10/Y OAI21X1_340/Y gnd vdd DFFPOSX1
XAOI21X1_55 INVX1_380/Y AOI21X1_55/B AOI21X1_55/C gnd AOI21X1_55/Y vdd AOI21X1
XINVX1_405 BUFX2_39/Y gnd INVX1_405/Y vdd INVX1
XOAI21X1_8 EN_request_put INVX1_17/Y INVX1_16/Y gnd OAI21X1_8/Y vdd OAI21X1
XFILL_25_1_0 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XBUFX2_58 BUFX2_58/A gnd BUFX2_58/Y vdd BUFX2
XFILL_5_2_0 gnd vdd FILL
XNAND2X1_121 AND2X2_4/Y INVX1_114/A gnd NAND2X1_121/Y vdd NAND2X1
XINVX1_369 BUFX2_28/Y gnd INVX1_369/Y vdd INVX1
XOAI21X1_548 INVX1_619/Y NAND2X1_522/Y OAI21X1_547/Y gnd OAI21X1_548/Y vdd OAI21X1
XDFFPOSX1_187 INVX1_38/A CLKBUF1_40/Y OAI21X1_285/Y gnd vdd DFFPOSX1
XAOI21X1_19 INVX1_128/Y AOI21X1_19/B AOI21X1_19/C gnd AOI21X1_19/Y vdd AOI21X1
XBUFX2_22 BUFX2_22/A gnd BUFX2_22/Y vdd BUFX2
XAOI22X1_96 AND2X2_18/B INVX1_321/Y INVX1_323/Y AOI22X1_96/D gnd AOI22X1_96/Y vdd
+ AOI22X1
XDFFPOSX1_151 INVX1_249/A CLKBUF1_35/Y OAI21X1_230/Y gnd vdd DFFPOSX1
XNAND2X1_82 AND2X2_1/Y INVX1_65/A gnd OAI21X1_68/B vdd NAND2X1
XOAI21X1_67 INVX1_62/Y INVX1_65/Y OAI21X1_67/C gnd OAI21X1_68/C vdd OAI21X1
XDFFPOSX1_85 NOR2X1_56/A CLKBUF1_14/Y NAND3X1_45/Y gnd vdd DFFPOSX1
XAOI22X1_153 NAND2X1_450/Y AND2X2_119/Y AOI22X1_153/C NOR2X1_202/Y gnd AOI22X1_153/Y
+ vdd AOI22X1
XINVX1_333 INVX1_333/A gnd INVX1_333/Y vdd INVX1
XOAI21X1_512 INVX1_577/Y OAI21X1_512/B OAI21X1_512/C gnd OAI21X1_512/Y vdd OAI21X1
XAOI22X1_60 AND2X2_8/B INVX1_195/Y NOR2X1_77/B AOI22X1_60/D gnd AOI22X1_60/Y vdd AOI22X1
XNAND2X1_46 AOI22X1_9/C NOR2X1_21/Y gnd OAI21X1_29/C vdd NAND2X1
XOAI21X1_31 INVX1_34/Y NOR2X1_21/Y NAND2X1_48/Y gnd OAI21X1_31/Y vdd OAI21X1
XDFFPOSX1_115 OR2X2_4/A CLKBUF1_45/Y OAI21X1_174/Y gnd vdd DFFPOSX1
XINVX1_297 AND2X2_72/B gnd INVX1_297/Y vdd INVX1
XDFFPOSX1_49 AND2X2_1/B CLKBUF1_21/Y NAND3X1_27/Y gnd vdd DFFPOSX1
XAOI22X1_117 NAND2X1_351/Y AND2X2_92/Y AOI22X1_117/C NOR2X1_148/Y gnd OAI21X1_358/C
+ vdd AOI22X1
XOAI21X1_476 INVX1_535/Y NAND2X1_456/Y OAI21X1_476/C gnd OAI21X1_476/Y vdd OAI21X1
XAOI22X1_24 INVX1_70/A INVX1_69/Y INVX1_71/Y AOI22X1_24/D gnd OAI21X1_76/B vdd AOI22X1
XDFFPOSX1_13 INVX1_9/A CLKBUF1_34/Y NAND2X1_39/Y gnd vdd DFFPOSX1
XNAND2X1_10 INVX1_511/A INVX1_469/A gnd NOR2X1_5/B vdd NAND2X1
XOAI21X1_440 INVX1_493/Y NAND2X1_423/Y OAI21X1_440/C gnd OAI21X1_440/Y vdd OAI21X1
XINVX1_261 AND2X2_64/B gnd INVX1_261/Y vdd INVX1
XNAND3X1_87 NOR2X1_100/Y NAND3X1_86/Y NAND3X1_87/C gnd NAND3X1_87/Y vdd NAND3X1
XNAND3X1_51 NOR2X1_61/Y NAND3X1_51/B NAND3X1_51/C gnd NAND3X1_51/Y vdd NAND3X1
XOAI21X1_404 INVX1_451/Y OAI21X1_404/B OAI21X1_404/C gnd OAI21X1_404/Y vdd OAI21X1
XINVX1_225 BUFX2_69/Y gnd INVX1_225/Y vdd INVX1
XNAND2X1_518 INVX1_76/A INVX1_608/Y gnd OAI21X1_543/B vdd NAND2X1
XINVX1_189 AND2X2_3/B gnd INVX1_189/Y vdd INVX1
XOAI21X1_368 INVX1_409/Y OAI21X1_368/B OAI21X1_367/Y gnd OAI21X1_368/Y vdd OAI21X1
XINVX1_71 BUFX2_42/Y gnd INVX1_71/Y vdd INVX1
XFILL_18_1 gnd vdd FILL
XNAND3X1_15 NOR2X1_20/Y OAI21X1_27/Y OR2X2_2/Y gnd NAND3X1_15/Y vdd NAND3X1
XNAND2X1_482 INVX1_560/A BUFX2_125/Y gnd NAND2X1_482/Y vdd NAND2X1
XAND2X2_120 BUFX2_63/Y INVX1_528/A gnd AND2X2_120/Y vdd AND2X2
XAND2X2_93 BUFX2_38/Y INVX1_402/A gnd AND2X2_93/Y vdd AND2X2
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_153 AND2X2_7/Y gnd INVX1_153/Y vdd INVX1
XOAI21X1_332 INVX1_367/Y OAI21X1_332/B OAI21X1_331/Y gnd OAI21X1_332/Y vdd OAI21X1
XNAND2X1_446 BUFX2_93/Y INVX1_520/A gnd NAND2X1_446/Y vdd NAND2X1
XAND2X2_57 INVX1_210/A INVX1_219/A gnd INVX1_209/A vdd AND2X2
XINVX1_117 BUFX2_28/Y gnd NOR2X1_52/B vdd INVX1
XOAI21X1_296 INVX1_325/Y NAND2X1_291/Y OAI21X1_296/C gnd OAI21X1_296/Y vdd OAI21X1
XNAND2X1_410 BUFX2_90/Y INVX1_471/Y gnd AOI22X1_138/D vdd NAND2X1
XAND2X2_21 AND2X2_21/A AND2X2_21/B gnd INVX1_624/A vdd AND2X2
XOAI21X1_260 INVX1_280/Y OAI21X1_260/B NAND3X1_89/A gnd AOI21X1_41/C vdd OAI21X1
XNOR2X1_96 gnd NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XNAND2X1_374 INVX1_422/A NAND2X1_373/Y gnd AOI22X1_125/A vdd NAND2X1
XFILL_11_1_1 gnd vdd FILL
XNOR2X1_60 INVX1_140/A INVX1_141/Y gnd NOR2X1_60/Y vdd NOR2X1
XINVX1_622 BUFX2_10/Y gnd INVX1_622/Y vdd INVX1
XOAI21X1_224 INVX1_242/Y AOI22X1_72/Y AOI22X1_73/Y gnd OAI21X1_224/Y vdd OAI21X1
XNAND2X1_338 BUFX2_38/Y INVX1_377/Y gnd OAI21X1_345/B vdd NAND2X1
XNAND3X1_170 INVX1_566/A INVX1_568/Y INVX1_569/Y gnd NAND3X1_170/Y vdd NAND3X1
XCLKBUF1_48 BUFX2_3/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XINVX1_586 INVX1_89/A gnd INVX1_586/Y vdd INVX1
XNOR2X1_24 OR2X2_4/A OR2X2_4/B gnd NOR2X1_24/Y vdd NOR2X1
XOAI21X1_188 INVX1_484/A NOR2X1_79/B INVX1_203/Y gnd OAI21X1_188/Y vdd OAI21X1
XNOR2X1_221 gnd INVX1_565/Y gnd NOR2X1_221/Y vdd NOR2X1
XNAND2X1_302 INVX1_357/A INVX1_352/A gnd NOR3X1_2/B vdd NAND2X1
XDFFPOSX1_368 AND2X2_21/A CLKBUF1_2/Y AOI21X1_90/Y gnd vdd DFFPOSX1
XNAND3X1_134 INVX1_440/A INVX1_442/Y INVX1_443/Y gnd NAND3X1_135/B vdd NAND3X1
XINVX1_550 INVX1_550/A gnd INVX1_550/Y vdd INVX1
XCLKBUF1_12 BUFX2_7/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XBUFX2_135 INVX1_16/A gnd RDY_request_put vdd BUFX2
XOAI21X1_152 BUFX2_48/Y INVX1_160/Y OAI21X1_152/C gnd NAND3X1_55/C vdd OAI21X1
XNOR2X1_185 gnd INVX1_481/Y gnd NOR2X1_185/Y vdd NOR2X1
XNAND2X1_266 INVX1_289/A NAND2X1_265/Y gnd AOI22X1_87/A vdd NAND2X1
XFILL_0_0_0 gnd vdd FILL
XDFFPOSX1_332 INVX1_562/A CLKBUF1_42/Y AOI21X1_81/Y gnd vdd DFFPOSX1
XINVX1_514 INVX1_395/A gnd INVX1_514/Y vdd INVX1
XFILL_18_1_1 gnd vdd FILL
XFILL_16_3_2 gnd vdd FILL
XXNOR2X1_59 AND2X2_7/Y INVX1_440/A gnd AOI21X1_64/B vdd XNOR2X1
XOAI21X1_116 INVX1_118/Y INVX1_121/Y AOI22X1_39/C gnd OAI21X1_116/Y vdd OAI21X1
XNOR2X1_149 gnd INVX1_397/Y gnd NOR2X1_149/Y vdd NOR2X1
XNAND2X1_230 INVX1_244/A INVX1_247/Y gnd AOI22X1_74/D vdd NAND2X1
XINVX1_478 INVX1_478/A gnd INVX1_478/Y vdd INVX1
XDFFPOSX1_296 INVX1_499/A CLKBUF1_23/Y AOI21X1_72/Y gnd vdd DFFPOSX1
XXNOR2X1_23 INVX1_190/A AND2X2_3/Y gnd XNOR2X1_23/Y vdd XNOR2X1
XNAND2X1_194 INVX1_484/A INVX1_205/A gnd OAI21X1_191/B vdd NAND2X1
XNOR2X1_113 gnd INVX1_313/Y gnd NAND3X1_99/A vdd NOR2X1
XDFFPOSX1_260 INVX1_436/A CLKBUF1_35/Y AOI21X1_63/Y gnd vdd DFFPOSX1
XINVX1_442 AND2X2_7/Y gnd INVX1_442/Y vdd INVX1
XBUFX2_95 BUFX2_96/A gnd BUFX2_95/Y vdd BUFX2
XNAND2X1_158 AND2X2_7/B BUFX2_49/Y gnd NAND2X1_159/B vdd NAND2X1
XDFFPOSX1_224 AND2X2_3/A CLKBUF1_10/Y AOI21X1_54/Y gnd vdd DFFPOSX1
XINVX1_406 INVX1_406/A gnd INVX1_406/Y vdd INVX1
XAOI21X1_56 INVX1_387/Y AOI21X1_56/B AOI21X1_56/C gnd AOI21X1_56/Y vdd AOI21X1
XFILL_7_0_0 gnd vdd FILL
XNAND2X1_122 INVX1_113/A INVX1_111/Y gnd OAI21X1_112/B vdd NAND2X1
XOAI21X1_9 INVX1_3/Y INVX1_15/Y OAI21X1_8/Y gnd OAI21X1_9/Y vdd OAI21X1
XFILL_25_1_1 gnd vdd FILL
XFILL_23_3_2 gnd vdd FILL
XBUFX2_59 BUFX2_58/A gnd BUFX2_59/Y vdd BUFX2
XFILL_5_2_1 gnd vdd FILL
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XOAI21X1_549 INVX1_616/Y OAI21X1_549/B NOR2X1_241/Y gnd AOI21X1_89/C vdd OAI21X1
XAOI21X1_20 INVX1_135/Y AOI21X1_20/B AOI21X1_20/C gnd AOI21X1_20/Y vdd AOI21X1
XDFFPOSX1_188 INVX1_310/A CLKBUF1_40/Y AOI21X1_45/Y gnd vdd DFFPOSX1
XBUFX2_23 BUFX2_22/A gnd INVX1_43/A vdd BUFX2
XNAND2X1_83 INVX1_64/A INVX1_62/Y gnd OAI21X1_69/B vdd NAND2X1
XAOI22X1_97 AOI22X1_97/A AND2X2_76/Y AOI22X1_97/C AOI22X1_97/D gnd AOI22X1_97/Y vdd
+ AOI22X1
XDFFPOSX1_152 INVX1_247/A CLKBUF1_35/Y AOI21X1_36/Y gnd vdd DFFPOSX1
XAOI22X1_154 INVX1_525/A INVX1_524/Y INVX1_526/Y NAND2X1_453/Y gnd AOI22X1_154/Y vdd
+ AOI22X1
XDFFPOSX1_86 AOI22X1_43/C CLKBUF1_2/Y OAI21X1_129/Y gnd vdd DFFPOSX1
XOAI21X1_68 INVX1_66/Y OAI21X1_68/B OAI21X1_68/C gnd OAI21X1_68/Y vdd OAI21X1
XBUFX2_1 CLK gnd BUFX2_1/Y vdd BUFX2
XOAI21X1_513 INVX1_574/Y OAI21X1_513/B NOR2X1_223/Y gnd AOI21X1_83/C vdd OAI21X1
XINVX1_334 INVX1_89/A gnd INVX1_334/Y vdd INVX1
XAOI22X1_61 AOI22X1_61/A AND2X2_55/Y AOI22X1_61/C NOR2X1_77/Y gnd AOI22X1_61/Y vdd
+ AOI22X1
XNAND2X1_47 OR2X2_3/B NOR2X1_21/Y gnd NAND2X1_47/Y vdd NAND2X1
XOAI21X1_32 INVX1_35/Y NOR2X1_21/Y NAND2X1_49/Y gnd OAI21X1_32/Y vdd OAI21X1
XDFFPOSX1_50 AOI22X1_25/C CLKBUF1_51/Y OAI21X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 INVX1_184/A CLKBUF1_49/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XAOI22X1_118 INVX1_399/A INVX1_398/Y INVX1_400/Y NAND2X1_354/Y gnd AOI22X1_118/Y vdd
+ AOI22X1
XINVX1_298 INVX1_479/A gnd INVX1_298/Y vdd INVX1
XOAI21X1_477 INVX1_532/Y OAI21X1_477/B NOR2X1_205/Y gnd AOI21X1_77/C vdd OAI21X1
XAOI22X1_25 NAND2X1_91/Y AND2X2_34/Y AOI22X1_25/C NOR2X1_38/Y gnd OAI21X1_76/C vdd
+ AOI22X1
XNAND2X1_11 INVX1_434/A INVX1_254/A gnd NOR2X1_6/A vdd NAND2X1
XDFFPOSX1_14 INVX1_10/A CLKBUF1_5/Y NAND2X1_40/Y gnd vdd DFFPOSX1
XOAI21X1_441 INVX1_490/Y OAI21X1_441/B NOR2X1_187/Y gnd AOI21X1_71/C vdd OAI21X1
XINVX1_262 AND2X2_66/B gnd INVX1_262/Y vdd INVX1
XNAND3X1_88 INVX1_279/A INVX1_281/Y INVX1_282/Y gnd NAND3X1_88/Y vdd NAND3X1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XNAND3X1_52 AND2X2_7/Y INVX1_155/Y INVX1_156/Y gnd NAND3X1_52/Y vdd NAND3X1
XOAI21X1_405 INVX1_448/Y NAND2X1_391/Y NOR2X1_169/Y gnd AOI21X1_65/C vdd OAI21X1
XNAND2X1_519 BUFX2_9/Y INVX1_611/Y gnd AOI22X1_178/D vdd NAND2X1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_190 INVX1_190/A gnd NOR2X1_75/B vdd INVX1
XOAI21X1_369 INVX1_406/Y NAND2X1_358/Y NOR2X1_151/Y gnd AOI21X1_59/C vdd OAI21X1
XAND2X2_121 BUFX2_65/Y INVX1_535/A gnd AND2X2_121/Y vdd AND2X2
XFILL_18_2 gnd vdd FILL
XNAND3X1_16 INVX1_28/A EN_response_get INVX1_27/A gnd OAI21X1_37/C vdd NAND3X1
XNAND2X1_483 INVX1_562/A NAND2X1_482/Y gnd AOI22X1_165/A vdd NAND2X1
XAND2X2_94 BUFX2_41/Y INVX1_409/A gnd AND2X2_94/Y vdd AND2X2
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_154 AND2X2_7/B gnd INVX1_154/Y vdd INVX1
XOAI21X1_333 INVX1_364/Y OAI21X1_333/B NOR2X1_133/Y gnd AOI21X1_53/C vdd OAI21X1
XNAND2X1_447 BUFX2_65/Y INVX1_517/Y gnd OAI21X1_465/B vdd NAND2X1
XAND2X2_58 INVX1_209/A INVX1_221/A gnd AND2X2_58/Y vdd AND2X2
XINVX1_118 AND2X2_42/A gnd INVX1_118/Y vdd INVX1
XOAI21X1_297 INVX1_322/Y NAND2X1_292/Y NOR2X1_115/Y gnd AOI21X1_47/C vdd OAI21X1
XNAND2X1_411 INVX1_469/A BUFX2_132/Y gnd NAND2X1_412/B vdd NAND2X1
XAND2X2_22 BUFX2_69/Y INVX1_5/Y gnd INVX1_27/A vdd AND2X2
XFILL_11_1_2 gnd vdd FILL
XOAI21X1_261 INVX1_284/Y AOI22X1_84/Y AOI22X1_85/Y gnd OAI21X1_261/Y vdd OAI21X1
XNOR2X1_97 NOR2X1_97/A INVX1_260/Y gnd NOR2X1_97/Y vdd NOR2X1
XNAND2X1_375 BUFX2_87/Y INVX1_429/A gnd OAI21X1_386/B vdd NAND2X1
XINVX1_623 INVX1_623/A gnd INVX1_623/Y vdd INVX1
XNOR2X1_61 gnd NOR2X1_61/B gnd NOR2X1_61/Y vdd NOR2X1
XOAI21X1_225 INVX1_244/A NOR2X1_92/B INVX1_245/Y gnd OAI21X1_226/C vdd OAI21X1
XNAND2X1_339 BUFX2_73/Y INVX1_380/Y gnd AOI22X1_112/D vdd NAND2X1
XCLKBUF1_49 BUFX2_5/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XNAND3X1_171 NOR2X1_221/Y NAND3X1_170/Y NAND3X1_171/C gnd NAND3X1_171/Y vdd NAND3X1
XINVX1_587 BUFX2_24/Y gnd INVX1_587/Y vdd INVX1
XOAI21X1_189 INVX1_204/A INVX1_202/Y OAI21X1_188/Y gnd NAND3X1_67/C vdd OAI21X1
XNOR2X1_25 OR2X2_5/A OR2X2_4/B gnd NOR2X1_25/Y vdd NOR2X1
XNAND2X1_303 INVX1_371/A INVX1_364/A gnd NOR3X1_2/C vdd NAND2X1
XNOR2X1_222 INVX1_567/A INVX1_568/Y gnd NOR2X1_222/Y vdd NOR2X1
XFILL_12_2_0 gnd vdd FILL
XDFFPOSX1_369 INVX1_623/A CLKBUF1_3/Y NAND3X1_187/Y gnd vdd DFFPOSX1
XNAND3X1_135 NOR2X1_167/Y NAND3X1_135/B OAI21X1_396/Y gnd NAND3X1_135/Y vdd NAND3X1
XCLKBUF1_13 BUFX2_6/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XINVX1_551 BUFX2_33/Y gnd INVX1_551/Y vdd INVX1
XBUFX2_136 OR2X2_2/B gnd RDY_response_get vdd BUFX2
XNOR2X1_186 INVX1_483/A INVX1_484/Y gnd NOR2X1_186/Y vdd NOR2X1
XOAI21X1_153 INVX1_160/Y INVX1_163/Y AOI22X1_51/C gnd OAI21X1_153/Y vdd OAI21X1
XNAND2X1_267 INVX1_324/A INVX1_317/A gnd NOR2X1_106/A vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
XDFFPOSX1_333 INVX1_560/A CLKBUF1_42/Y NAND3X1_169/Y gnd vdd DFFPOSX1
XBUFX2_100 BUFX2_98/A gnd BUFX2_100/Y vdd BUFX2
XINVX1_515 INVX1_515/A gnd INVX1_515/Y vdd INVX1
XFILL_18_1_2 gnd vdd FILL
XXNOR2X1_60 AND2X2_8/Y BUFX2_113/Y gnd AOI21X1_65/B vdd XNOR2X1
XNAND2X1_231 INVX1_245/A BUFX2_15/Y gnd NAND2X1_231/Y vdd NAND2X1
XOAI21X1_117 INVX1_122/Y OAI21X1_117/B OAI21X1_116/Y gnd DFFPOSX1_78/D vdd OAI21X1
XNOR2X1_150 INVX1_399/A INVX1_400/Y gnd NOR2X1_150/Y vdd NOR2X1
XDFFPOSX1_297 INVX1_497/A CLKBUF1_23/Y NAND3X1_151/Y gnd vdd DFFPOSX1
XINVX1_479 INVX1_479/A gnd INVX1_479/Y vdd INVX1
XXNOR2X1_24 INVX1_197/A AND2X2_8/Y gnd AOI21X1_29/B vdd XNOR2X1
XNAND2X1_195 INVX1_204/A INVX1_202/Y gnd NAND2X1_195/Y vdd NAND2X1
XNOR2X1_114 AND2X2_12/B INVX1_316/Y gnd AOI22X1_95/D vdd NOR2X1
XDFFPOSX1_261 INVX1_434/A CLKBUF1_37/Y NAND3X1_133/Y gnd vdd DFFPOSX1
XINVX1_443 AND2X2_7/A gnd INVX1_443/Y vdd INVX1
XFILL_19_2_0 gnd vdd FILL
XBUFX2_96 BUFX2_96/A gnd BUFX2_96/Y vdd BUFX2
XNAND2X1_159 INVX1_156/A NAND2X1_159/B gnd AOI22X1_49/A vdd NAND2X1
XDFFPOSX1_225 INVX1_371/A CLKBUF1_33/Y NAND3X1_115/Y gnd vdd DFFPOSX1
XINVX1_407 AND2X2_5/Y gnd INVX1_407/Y vdd INVX1
XAOI21X1_57 INVX1_394/Y AOI21X1_57/B AOI21X1_57/C gnd AOI21X1_57/Y vdd AOI21X1
XFILL_25_1_2 gnd vdd FILL
XBUFX2_60 BUFX2_58/A gnd BUFX2_60/Y vdd BUFX2
XFILL_5_2_2 gnd vdd FILL
XNAND2X1_123 AND2X2_4/Y INVX1_114/Y gnd AOI22X1_36/D vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
XAOI21X1_21 INVX1_142/Y XNOR2X1_16/Y AOI21X1_21/C gnd AOI21X1_21/Y vdd AOI21X1
XDFFPOSX1_1 NOR2X1_10/A CLKBUF1_9/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XDFFPOSX1_189 INVX1_308/A CLKBUF1_40/Y NAND3X1_97/Y gnd vdd DFFPOSX1
XINVX1_371 INVX1_371/A gnd INVX1_371/Y vdd INVX1
XOAI21X1_550 INVX1_620/Y OAI21X1_550/B OAI21X1_550/C gnd OAI21X1_550/Y vdd OAI21X1
XBUFX2_24 BUFX2_22/A gnd BUFX2_24/Y vdd BUFX2
XOAI21X1_69 INVX1_63/Y OAI21X1_69/B NOR2X1_35/Y gnd AOI21X1_10/C vdd OAI21X1
XNAND2X1_84 AND2X2_1/Y INVX1_65/Y gnd NAND2X1_84/Y vdd NAND2X1
XAOI22X1_98 AND2X2_21/B INVX1_328/Y INVX1_330/Y AOI22X1_98/D gnd AOI22X1_98/Y vdd
+ AOI22X1
XDFFPOSX1_153 INVX1_245/A CLKBUF1_35/Y NAND3X1_79/Y gnd vdd DFFPOSX1
XAOI22X1_155 NAND2X1_455/Y AND2X2_120/Y AOI22X1_155/C NOR2X1_204/Y gnd AOI22X1_155/Y
+ vdd AOI22X1
XDFFPOSX1_87 INVX1_129/A CLKBUF1_2/Y DFFPOSX1_87/D gnd vdd DFFPOSX1
XOAI21X1_514 INVX1_578/Y AOI22X1_168/Y AOI22X1_169/Y gnd OAI21X1_514/Y vdd OAI21X1
XINVX1_335 BUFX2_22/Y gnd INVX1_335/Y vdd INVX1
XBUFX2_2 CLK gnd BUFX2_2/Y vdd BUFX2
XAOI22X1_62 AND2X2_10/B INVX1_202/Y NOR2X1_79/B AOI22X1_62/D gnd AOI22X1_62/Y vdd
+ AOI22X1
XOAI21X1_33 INVX1_36/Y NOR2X1_21/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XNAND2X1_48 OR2X2_4/A NOR2X1_21/Y gnd NAND2X1_48/Y vdd NAND2X1
XFILL_26_2_0 gnd vdd FILL
XDFFPOSX1_51 INVX1_74/A CLKBUF1_26/Y OAI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 NOR2X1_73/A CLKBUF1_6/Y NAND3X1_61/Y gnd vdd DFFPOSX1
XFILL_6_3_0 gnd vdd FILL
XAOI22X1_119 NAND2X1_356/Y AND2X2_93/Y OAI21X1_361/C NOR2X1_150/Y gnd AOI22X1_119/Y
+ vdd AOI22X1
XOAI21X1_478 INVX1_536/Y OAI21X1_478/B OAI21X1_478/C gnd OAI21X1_478/Y vdd OAI21X1
XINVX1_299 BUFX2_33/Y gnd INVX1_299/Y vdd INVX1
XNAND2X1_12 INVX1_553/A INVX1_518/A gnd NOR2X1_6/B vdd NAND2X1
XAOI22X1_26 INVX1_77/A INVX1_76/Y INVX1_78/Y AOI22X1_26/D gnd OAI21X1_82/B vdd AOI22X1
XDFFPOSX1_15 INVX1_11/A CLKBUF1_34/Y NAND2X1_41/Y gnd vdd DFFPOSX1
XOAI21X1_442 INVX1_494/Y OAI21X1_442/B AOI22X1_145/Y gnd OAI21X1_442/Y vdd OAI21X1
XINVX1_263 AND2X2_65/B gnd INVX1_263/Y vdd INVX1
XNAND3X1_89 NAND3X1_89/A NAND3X1_88/Y NAND3X1_89/C gnd NAND3X1_89/Y vdd NAND3X1
XOAI21X1_406 INVX1_452/Y OAI21X1_406/B OAI21X1_406/C gnd OAI21X1_406/Y vdd OAI21X1
XINVX1_227 AND2X2_60/B gnd INVX1_227/Y vdd INVX1
XNAND3X1_53 NOR2X1_63/Y NAND3X1_52/Y NAND3X1_53/C gnd NAND3X1_53/Y vdd NAND3X1
XNAND2X1_520 INVX1_609/A INVX1_76/A gnd NAND2X1_520/Y vdd NAND2X1
XNAND2X1_1 INVX1_336/A INVX1_44/A gnd NOR2X1_1/A vdd NAND2X1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_191 INVX1_191/A gnd INVX1_191/Y vdd INVX1
XOAI21X1_370 INVX1_410/Y OAI21X1_370/B AOI22X1_121/Y gnd OAI21X1_370/Y vdd OAI21X1
XAND2X2_122 BUFX2_66/Y INVX1_542/A gnd AND2X2_122/Y vdd AND2X2
XFILL_18_3 gnd vdd FILL
XNAND2X1_484 INVX1_566/A AND2X2_16/A gnd NAND2X1_484/Y vdd NAND2X1
XNAND3X1_17 NAND3X1_17/A AND2X2_26/Y AOI21X1_6/Y gnd INVX1_5/A vdd NAND3X1
XAND2X2_95 BUFX2_38/Y INVX1_416/A gnd AND2X2_95/Y vdd AND2X2
XINVX1_155 BUFX2_49/Y gnd INVX1_155/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XOAI21X1_334 INVX1_368/Y AOI22X1_108/Y OAI21X1_334/C gnd OAI21X1_334/Y vdd OAI21X1
XNAND2X1_448 BUFX2_93/Y INVX1_520/Y gnd NAND2X1_448/Y vdd NAND2X1
XAND2X2_59 BUFX2_55/Y AND2X2_59/B gnd AND2X2_59/Y vdd AND2X2
XINVX1_119 NOR2X1_53/A gnd INVX1_119/Y vdd INVX1
XOAI21X1_298 INVX1_326/Y AOI22X1_96/Y AOI22X1_97/Y gnd OAI21X1_298/Y vdd OAI21X1
XNAND2X1_412 INVX1_471/A NAND2X1_412/B gnd NAND2X1_412/Y vdd NAND2X1
XAND2X2_23 OR2X2_1/A AND2X2_23/B gnd AOI21X1_1/A vdd AND2X2
XNOR2X1_98 gnd INVX1_264/Y gnd NOR2X1_98/Y vdd NOR2X1
XOAI21X1_262 INVX1_575/A INVX1_288/Y INVX1_287/Y gnd OAI21X1_263/C vdd OAI21X1
.ends

